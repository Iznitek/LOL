MPQ    ��    h�  h                                                                                 9I=Nʂbd�X7n'��
x�{tLGY����7�E�a�u�S�k�\��W��޷l�dJE�6���U}x�]������'�]dB�#Ŏc��=|��[����<�Y�W�Z�Ϳs%��Qmz�I�!ck�A>ԭ6�x�)_Z��$;��ae�����p4;q_��}�N��5�����*N��f0�kR�3 >k�[c��H�3�-����K/�)�E�!�U�Cڴ
Yx�i�zkS��dl�W�R�9R3�0�rHg$�7�F����/ׯ�f3Iu>%��:��8�C�����I��k�F�#A!�����\�����G�h�bw�~�<w�]/�N�:��p�� �Ɉ��m����\��]r���"���+��=w���!}<xҐ����B¾�Z|�S*��s���H;ƍfy�c[����-O��qy���S�|��B���J(�EA�V��l_�l���	��&_=��Lλؑ!�&�U��hK6d����|����s8�kC�˚\#���cZl7ډ�-')�U��B���T��/������@ܕ���7�+�e���3��us��{ �˒��-�g�@Se�<�2���ɉ��kS���lgv1*2}1ba�i���Rķt��ŀ#,`�h��t��J��
J�m���2�b?�c�Hy�M#�@k&�ߣ�ygX�/n�/W��E�a��aYs��{�~N�,
��9��~l���Uq�������ݖ0oT{(�{��E�.�k:!V�ve=%��C��Y{����/���u��,[^�9��1���S��%&����ߍZ�.�5v�g��]IW��'��X@��G�l����.�"��x���N�������tS�`յ $����4��o�3Tw�t�	��+�te�b����H@���?*`n!,���?0�Uj��}u:f���g�������o&�+d�b���V�-+ڇ ��.����c���)w���ẁ��d���͒&e����_��V�Jh�P�Z*�l����U�˨�m��o��
���?��3�2L��!~< �e��Sx�ǡt��������V���$��H.�Vp�jI�Q�=pj7�#B�u����hXd��:�����{@�-����(GV�����(BV�
���<��-5!=���P�c�LY��I���������,���B�Ĭq�^*a���'�5���k<x�����Yj>(a�}��{7�qr5w�m�T]��{ϗ��c�Q�	(�~�$��œ��Zq�G=iJ� �QM�^j ,�0�I�S��?B���́ψ������C?��Ȕ�U����m$�J�ц�@ 5�`�S�&#��V��ֆ �6�n�k�gI\�A���c��6 X��#{�!i轿&�w��Y̿��>h9-MW-�׵q.]-MV=Ϭ�a".Jp^�p�l+��yc��ō���-�����C�d�!	���z;�A7����|;|�ܳ�ۈOm��1�0+��Sf@��'/#V�"���2��	�Oz 6l�����@n;5�p�����Q�Ь�'�%���pW�!����C���	 �XNo�Y'?��	�sޜ���w,�!Ģe�����]B���y�w�uk��8�ۊ�/��iu�C�}�y�K�󂦰�z"O�y�m�l栾�zF~��O�G�I�2��� �t6H��!r\�&��=�OQ�Ȝ�W��⪫�=�����R��J5���M�^�`�?�\�X����?N���o_��ǖ��~R�0U�hP�	t���/�ЙL�ڨ��[��4�eq���y/��2���Z�� �m�ϋ��<�N�%�ǃ8���4����L9���yAg��*�>nei�*0�WY��3� �:��PǑ4+$�Hc���ÏJ��5�e�q2_P�Z'e�/-=E���c�M���'�	�1xpJo{8�=Y�s{Q�I$s�+'F+����1����7-H��-�ia��u)�xR{�gh���g�=����͟�2q�en�	�;Ɵ�s2��:�Z�|t��6'S�<1��H))��K@��I��9��	<<>�Vo�_г�A��'�E�P��?���j��"�DD
��FAL6�0���.
K�e��s�P�о>��+�E�	��|�/K#��*���Y��F���(<}�J7�z�Ӏ̬�1(�J]���uؔ�틉���f#�He�n�`R��J,#6�Xf�,x�ܠ�6�E���0c��u�ά/�c
��2W�K����"~��m �P���rkM�|cŗogJ5�~��r�����F�A���]�/�p�8�l�m��-���#����Ӑ�f���b���W�/�q��+��dU\�
�ح�%�/�%º�lT?٭[��q���k}�˛����Yn5N��H��D�����c���O�XC��#Z#~��c:���i�"踿F����4�����w�u�N���u��p��jZ�Ҧ�BU ��s��G���|�� p.����{�i�Ua�2����Vv+�^�zA�q��hZ/�)Uy�n�����w�T��˘M��5�B���~y��-p��KJ��J���+�4�cM� A�C�9��[a��.t��V��!ɷ�woS��Q{KJ���h`�`xOzi��h"%ީǵL_V�V6����
#b��[K�e�p)��o`8̆�;;'˒��uP�k3�Zz�������؏zG��)��Ԝ�8�Z�'w�<���\�J'5�d�S��Q�.����'ټ����3;Q��F��+���	����u����4�އՙ�����z�%gmal��2]�	��@����ܛ�]ÅՆxw�q���f��'�9���UmZ:����"|��k������j��@��y����rq�@�f+8?�C�� ���æl�GT�j��J�F5?}���~O����rޜ����H���(��dEۛ~X+ 'T�H��g0�Ǚ�l�<�ʎ���JJu�yZ'�C�M�J�?�^��DJ=���ݯ��xp����'�z��նy�}ew�����R��dH0�x,ҵÛ�xyK@�q_�ړ��f�$�"+�0QVr2�h
��ّ��FD����E�>P��|]j�6�oˊRWB��^��=���[x֓(X����{0M�b�s��Q��I7}3k��>ԋ�y�)Z���8�O���a�Ʋ�s��p��_��F����5�Vf�F۪*	M�fK<C�3�^�k�{͍Dh�.�E�'��K���)�^�!��C��5E����fU�����WX�9V�̫"�HB��7R��2B�*�;�%�1�@A>@|`�U�Z�C�ƥ.N ��ߴ^ݹ#���}���y��eI�!K��t��yZwNx'/��P���� { }A��y�m�bx���Kڄ�8=�FŦ�����6}׽됮�8���?�7 �nŰ�������ﮂ������O���4���n[�|3�f��;8煼$E��E�	n?_�ڦ�NCW�A�6�F�����;����U�+�hz��d�w��7}y���2��"��u+%���Z)���R�'�U	߭_n�#�T�.	�
"&�+l�=�F���T7�b� �z�N��u��VE���IT-A/W@N <3MM�a�ۉ04��ƣp<vl�2d�a����*���/����o,ۭ5�]��� ����m	6��b�	Ȟcl�M��kᜣ�ZsaX*�9��a��L�a���Y�7{s�N�v
1U09 ��2����*q��;����o�rc�p[E����
�:�r�v��R%V*�C� �{����X��{o���U[��9k�1�&�S~��&07�Q�U'篐�UgK�GIr��ܢu�XMIGM�W����)�4��M�T�N���.	o��S�����P���;�O�3�
�m�	y�+�G���B;�z����ևO�>?�3S!G\3��s0���M�}�{��V)����G^&�a�ݤ��1�M+�E�t�x��Qm���Y��*��5ƕ�8��W���\&����_@��z�#\L����=A��NU�m��hz�o<si±�l�} ��&����#;�eUԬx�gt5��㪗���8�]���������j�O�8�7��{�04�6.d
 ��s$϶�
-*����GcK[�����C�ȅ�Kͣ�g �h�G=>ԸP�d�L�%����51\������,�w�B%}�q�*�(]��<���I<��N�����Är}�v���%r�v���q ]e��{��򳞒�/��(��$;#̓f�5qҫqi��,$�^���n*RI��|�K�������V"�����z~��c�pU�����Jϝ��zw5M�KS�SQ����'�� t=���k�:+Iw@A��cgu-6;+���!dvi���!w^�Y��V��h��Wh����s-H�(�D�"�͕^*�F=|+x��c"�J�(�#�(�m�`�CBst!$��M�W;���x���(�ע$�p�BO(1�1���YH�@�v�/^U[���O��N��
�c6����4�ko;p���10.�L?ɬ�K������;�l���_�~3*�x�g�S�Eog�'��	���ΎR�_\�:ev!���~���4�K��4Y��e+����uB�G�x�����=�_ѕ����64�G�4�,�z�{ש� �Gfǵ����tDt��������a c=7�L��W��Z�f���X4�<�>�h{��#BM[2�`��h\Up��re�Zw��T��â�ז�O�RRo�cbmZ�׵۹*�Lir&ȯ��oAM ��Ԝ/S���Ȩ����mL��s�É?A%|��8�t45y�Y߄�'v�y��3��n���*�8�Y�Z/�{e���nk�O�R$)���j	5��?���۬e����MRZ�q�J�Ed��c�7ʛ��K��l5,
��r�{�ԣY��Q,X�sp	+Ff@aLp�1��sϒ�m���Wi|*�����x-�g���ũ�=�A��(2,��nϔ.�7�;��6sm�K��z9�w�=���S���1�	w)���K�`49�ԭP	7qK��CC_��A�0"��O=P�j�?�Ґ���4�"
���
~��F\����b��c�K�5�����ˉԼ`�\+?��	��?$ t#^�m�	���e�����F`7�{�����(�Ճ���usB���"�������q}�۸���#q��Oq�'��7L_��-�s٫��UJ��j������W"G��e�2���xjK �ܯ�,z�Mdk)Œ1�g�1�9(��� �� �!�����]���p��Zl��۪�⹟Fɱ;t,�k�4�͝�b�zi�R�}/>m��nJ��\`�$؈��j�%]�l���D?40P��?+�2W�}SF��\��Ӕ�^5��H��D�g9�lpK��)C�Ӷ��<�~���:H��i�@}���)���4PѬ�s>�����]WOut���j��߈�U�� s���2��B�� k}g�MN�6�i�F)ast�����V�����A���ó��Yy1�H�V�f�%w����fJ�M���i�8B��$~��-��K�H]�ؿ@�f���C����sci�A�59E�[<��.�$��ݒ��ӷ��o'Q�(��GD�`a�OTA�w[�%$��R/��VQb�C��#=	�[��F����jq����|;��Î����3�"�KH�r�H�J�i�'G@�])U��O�F8d�'�`���"V�E�T��Bh�E.:�ݢ�����73<�n�|�ƨ��x���ą����r�
���,�;���u#rg�=@zP�xF�_��od�i�]�7�Ձ�Cwv#.�,���#��
����u���cm�O��a|����}&���B��T��ؠ%r�Сa��?/���� c���@lwk2��vׅ�;5�2<����O5���Z޷���z��eR���Ev�NX&T�T�\ß��1��
&W������<J� �yU&9������yv@D�N$��D����2���h'��zh�*���ye�H���#��ǿ�d20�T,-�̛�8Oyf��q�=��⤚fJ�"ưDQQҿ��C�W$��[U��՘���y��C;�]e����U�R��y=�=r��[SOޓc������v&YTus�+�Q�J,I���k��h>JU����)Ue�Ǔ�����a�)���e�p�F�_�,���x�5��\ס�r*�äff_4�T�3֟�kA�G�((��)6�܂�K���)�i!���C�l.��ҟ�aw��WL&98zi�&�mH27�~ɕ���%���_0~X>[�3���a�SC'���r������#�4�5wH�y��sRBa����t�3w�Z1/}	����f� X�k#�m]��Z��gX"�?nBXY��!�W�����h}r#����v��A��zHى���i�K�]C��x��܂��x�O@6��W}��|�;���ԕ��p5Ew4m�N_Vi��	���\ax���i���%�
�U#҉hu�d?1���a��K��a"y�P�Qm�Z�:���� '�9��hϞ�>h�T�x�廚�fA��I����7M*���|��i;�ui�c�1�c�*-�n@I�<�����2�Kq�a�ԣK,�v��g2��Va�������	����,V��8'����@��m��L35b����~�Mx1k�&�\i��%ƴ�D�Ns�a��7Yi�b{N�;N%�
���9��4T�t�q�s���a����oʉrͱnME��5�Rc:���v��%сC�g`{���e����C<[��K9-*O1y�nSY��&k8���h)P�;��$7gVI�H��c�X���G�1w�*�$-�a}��2N�����f^J�S2ǋ�6Y~��Ī��3�(����	���+l:��ؐ��*铺i���*?�'�!bǺ����0aq�N��}������x�]�r��&� �X���5+P0��~��0��=��.k��*��,��N�O�F�?��$_ql	BTq�>���������U4/ �co@o���l��!�U�(!����v��e� �x�'3t�G��eB]��:����۩H��pj��3f7@����9��##�d��%�N����V�-�ࠥS�G�`[�n���^�#� '����qۣa�=�A�P腅Lf-��0��P�.��G�Ԅ��R("B�U^q��Zǝp�0O<;
�ѿH���E^ȇ}�-�푚rx����
�]�gZ{�1��Y��@�(�b�$�䲓!��q�/i@��Y^��Q	DyI�͆��7�W�k�GW�0�\g��[���}�U�c�#3PJ��+��Ԗ5�{VSh����� W �$[k��2I��A�� cBm�6v��Y�!_$��[�w1�Y ��4	Zh�R�W�������-C(�b܎"�q?^E�$���+S��c]F����#�OԻaFC���!?�uȎa;���ʲR�ұ��˗�O��1�@��\4@��/�t�X��x(��%����6���|�F��;��~�̡԰G�=�Z��w���ަ��Х��h��G�N!o�'�U�	���|�G-V7�$ecu��\��Y��c�̽��C�@{@=�u݈K�s������gsѰj�o���"�8�gI%z|�ũ��]G�����	�(��t,��םqߜa�=�@`����WO�r�!��s����V�C̽�^��M�%a`��Z\�ů˂���u�ǡ�(��}ǫR���^�z��V�p�j�E8L�)Ȋ���Â��d���;/��/�[����Pm�9�NI���̆%�8�<�4g����B�y7�Z���0n�y *f�&Y�����WN�Z�S�j�B$�Yt�E������k�we��k
Z��,�e;E߂}ca���20��?��'3�&�q{�(�Y��Q���sK�F��t�P1�vZ���2�L��i���k�ox�fg�V!�D��=� �߃��2�URn�5����;|'�s�p��p1p�rhK�왯SP��1��)��K��o���o�5	2�ԧ8�_F�A̧��;�P��?�"�%d~B���=l
9�Fw���&����K&& ���~��t&��0�+�PW	����h#9� �D�� �Z��t�3��7H��	�4���(��2�Ou��k��y�P�6���V?�����#��ۅ�Ҙ"�����������&���VY�"7Y��>w��DWbQR~��M����� ��3�g��M�yGōqg 1��Y�������9���8�9Pu]3�p�r�lq�S�e�������&�F���<b:_ϑMO�/��3�c��ɚ��\��h�c�|ǥY�%�9ϝ���?�҄�^-��M�p}Ύu�7����5�:FH��DX5,�'闑���NJ0��?�~�C�:���i��ظ��}-�4˯��N̔��^���u�@`&�jБ�����U��sze�mn/�� f�HG�]��-�i��Ea��2�t�	V�	�j�A��?�-�*ByL*�|��A8bw9I���M��>��]�BJX~�+S-f��KŢ܃U��=����Y�=�rc�#�A�G�9���[�,.�Ĕ�L�$�7��m�jo�` Q�%����`<�O��l�n�%�T�kw_�m#VlJ���v#d�[�@���}�e���<>;�b��aF��3z���ι�؏�UuG�gZ)!��8?�'�,��+v��@����<�U�.1��R��rA^3w�`����/=�CQ��	��}����mu"���y�����p�:g#:5����
���0J�D�RV�]L̖�|��w�Jz�筘�����V<���P5��m�Ѐ�T�|R��h��4]��>�/�y���r�I9�\�G?���vI@�$�l���\����Ĥ5uǭ�p�O�4��������v��E8�@����[E�6X!��Ti�W�Z�6�L�������P�1#9J��TyPE���A��S���wDsW�w�<�6���l�q?'W>�z#d��y�em�q��q2�����0��,�>֛T�y��oqU������fW�"a��QLR��oG�����!:�d��4���Ѐ�ޒ$]`H��% �R�鎔�=�E$[.�6���F�*n�q<A��_sV�BQ��!I-��k��$>����I��)PF���'l�Ya���iL�p���_:����5��o���*Zf��Tu��3� �k|p���+P�$�*��twK`K)�7!kpCkx�����:�$\���u�{W��'9S��̡��H��67���hդ �y��/9��>v���K<�6CbQ�d��ଚ�l�#r��P����N_k��Q��3�-�oC�w]{/8W!��Ť�1X 3�U^��m�w������F�sI�Ŝ����?�P�:}���Ӱ�Sk�����٤[��)��8�>bւ4͙��|�O��Q�F��ǥ|)�3�u����D�E�̽��_�0���w�<j)�i]��Ed&U��lhp��d�
cӭf���_��A��+)���W�Z=lU����':>q�#_��Y�Ty���u��6�s��{ޔ7�Y�����Ƅ�u�f����C*�-w=@D��<��k��'͉f�������&<(v��2N)�a�[������8_���,�$����O-��ۂ�m�7����bpa����M��k��ǣI}�8�� "L@�ǃ	��aӦ�Y���{)�"N@QT
g��92n׏��/k�q�|�1!�njo�U�L��E����M�:Rnv��&%L��Cj��{W�� L����잘�[C��9H	A1�S4��&��s�]�K,�F�8g���I�ܘpkXѦ�GÉʥ�m�����/�<0rN�Z���%LSm*e��#�������3���ō�	�O+GM���;���鎣����?[;�!}RJ��i0</��A}F����� ��!��-e'&.���U�睞+�������/0�tO-�F��I���+��b@�։Uϒ�)���n�_����L�Y�F��h�����V�U���^�o�&�'C��<�2��;q˲["�+�e�M'x��t�&�� H��\ӹSQyۄ'�!�jer�.�7��憐��>02d AM�)���,b-`.�
�(G���)b�y�f�{"%��S��'�=tϏP��^Lj�.�z��k�	�����܆��DB[N�q�"*r��Xg6�+�|<��񸬀"�
�W�+�}��HH�r3Z����/][D{`{?�Aie(�B$��y�܌�q�i�����1^w��}I�:�PD>�(A� �����7)��X�ݙ"UzϘ�~j,JEÎ�O^5C9SC>�R:�]�� Z��akFv~I���A���c�;6�1���!Z�T�7�|w�iTYP[�\�h��W��d�B�->��Ͻ��"_5m^`3�P+.k�c�*��^)��^N�EC��!Z��Cx�;`, O���M*���P�&��O��1"8�O�@e޶/Գw����
r-�_U��H�6�{��*�J!-4;�*��g3�B�.����2�>�ƚ��-��c���������I��o6'p�2	/���ج?҄e�ʁ��y�SaҪ��"M��*����@<��ux['�n��\d�����˺���m���֬���z׫���G��I%�Cz�t��c�c����E=m鋵�pCW�3+�ܱf�4�2+��=��:M�9`�t�\,��=�y��):�J���X
j�X^�R�L��Y��#]��+[޹`l#L_f�eP��e�6���V/	n��8Q�^omB'@�)����y�%�ei8�$k4��ƣ�d��]�y�O.���qn2�*�"Y�Z�1j8�
�����$/� y�����e���p�"ZX�L����EZ�:c<��m����wH"|,�#�{i��Y2�Q"Վs&%�F���Q�1��]�H�����i����敂x�u�g;@��I�=}�4��zJ2��nn�Az�e;W��s�_Y���m��G�NS�1B)���K�<$�؀�
�	-;ڧgL�_3OA�>�Զ$lP���??�ȝ�jy��U}0
�0F�r�����z-)Ka6��D�)��4���+�	�*#����2��n���J�Q�7�O$)Ŭ�V?(�K!m�/u����|,��G'�MK�'؅���%�Kl#�0����\"��egi���A�١�#��w�]s��4���Q�W�.`��h��n× \T���VM���ň�g[rɺ����ÿ\�	���׍��t�G]Μ�p�?>l�R�� ������1���!� �C8�b�c͑H�^/�{��T�ɵ�\VY�>�p���g%��靜5Y?���;�h�}I����%�
h5�H���D�"��H��i���i��b#~1�d:~+�i�^3Ѽ�8Q��
$54F���)�{�&������u�h�G�j�@ �u�U� �sU����xq a{f�
-��g�i��ai}%�O�NV'��/��A��y�[�Z�yg�f>\��wt�T՜}M�Y�"�Bo�~�rt-���K�l�N
*������Z����c~��A�y�9^[�.%����Ln�����Do��Q�BP�=�-`p�O�{쭭�%��Ƽ��^�V�R?9�#��m[�d�A�`�`�I̗�;X�T�Tz�M�3��b+�¨�B񇴂��bG�n�)9��E!8m�'(�����;|H�u�����.L�hݘ>c�M�T3��&���x���]��B:��2|�x�<PIP�8|.�q&��k�~g~V��-�)W�Uh%�5��c�]��w��w,��ʢ��A� $IӰO�p�m+9	��g|�z��#ٽ�:��8*��
Q�N�IrB�y�We�?�O�1���*�-lm��7����5�I���O����<����-a�p�k�.t�5K4E�]7X�T����$0�gR�� �»�ě�lg�JxyK��T�[�{=���.D����R̤�q_#A��{r'��;zކ��ʅ�e�G����1�\�5�o0��5,�ߛ�y�ŧq��ړ�خf��^"��4QG������.�<�j�u	���@�y
][�����xR�#g���B=h�~[	/ߓ�i���Pflr
�sM�Qٚ�I�O-kk�P>�D���)KG!�I��'��a�O;��Rzp�һ_u/���
5�Z��W]�*:$f�[���-3��rk���^O�D��8��K[�)jN!�VCF���5z���W���1-W��9n"@�yHӿ?7���>	S�6�-��>�	r�D��*C�ܴ��ʸۤ�oc.#-��k�d�o�8)���3+�΃��jw_/���b�\�x i���amT��V��Rڵ?��Y������q�}�N��,献���Fb%ٿV[�_� �@��yKȂ��ȱ���O�\�eU�鿭�|�n��Pfa�69sE�d���_攲���ӝ�^5�D�j�cUY�hksld���h�����W�!�X˞�aZؽn���+'�b%���t�T�m�ЛO���K#s�v.7�~�Q�(Ɵ?:u_<g��s��~J!-F�@?"<D\[����K��WW�l�v��2黫a�A�;(��`��1a�,L�%��Η�c��v��m�����b+=���M�Rk�5����:�������  a��Y_ܤ{�N{��
p�9
yo��E��\+q���m��IF?o@���9E������:�$v�ͬ%ǐ+CEU'{�WLݛ�P���D���[���9c�1onVS�&��/�"r%F����SZg|!�I��<���X���G�R�`��ӿ��M!N�/B��7m ԝS����lb���x�`��3@Z�M[	�c�+"�e�N��KZ3鉬��`�?o!��ᴃ��0�ĸK}�|L��r�.u^��#&#�=�NQ���&�+�X�E3���k������[�dMW�S{=t_��#�|�z��ط_'�<��
�t@���W��z_���3Uj8�Y�toM�����W"��v�ˍ�9��e&�Hx�5tF&����V�񞿹����_\"�B�Bj�<��)܄7���a&�Y]`d{A�dZ�g�-�E��_6Gt�{��b�֔⑅�=��`���t=}oP�'4L�F��5(�������³�Ќ����B�fpq�Nb��5�~)�F��<~��a��E���Z}�����r���ٜ�]�@{;�OH ��(��$L� ���q#�i6����h�^V�G?�/I���p�����;���5֐�+v��4��Uu'j���(J �&��5�pS����7���Ԋ �|���?kDI�o`Av¨c��:6�dg�%K!U������w��GY8���*��h���W|�݄�-9z��m�"^{_��W
+	��c�s�������h�qH|Cs_�!u�����;;e������~��/A����OY�E1=5w���2@@/D�� P���_���;��6ؗ�奛N���;!�]�剰=���y�x�)���*����/3��I���DN�ox¿'+k�	J|��r���v<eGRF���J�;#�e�_=*N��z���z�w3�uNۈi��iT�n����%�e9�����U�z�4���ӵGw���as�^-Yt"�S��I����=�ϵ�L W����x�橮���������M,m�`��\f�n��*������a��3F떓)R#�B�TX�~���76�{�vL��'�@7� (��ט��+�/dJ-�џ���m�iӋM��:GN%Mڐ8�,�4띣�W@�x��y-ݭ��.�nQ
*�w�Y�s����b�Ї�-{$�굠�`j�6���[�e�)���Z�Ж���Eթ�c�⛨�n�u-��`ܫt{$0�YM�^Q�Cusc�F�Xri1��|ϣ:����iͬ�aO�x�^�gT?�z�=x���9Y�2]�On �7��;2/�so�զ���h�z䢌�S�)d1*s)-Kt{n��ڥrh	(�[�__��A�A�1�UP��?z₝[�ht⾷��
�{�F�,���UK�fF��������q%�+p�	:�1�#���β6���@o��7�=<?�=�	��(\6��
�uD��wͪ�/(~�7B;�L����#"k� {���c�H�"����$����q��Θ�S���Ĺ��FWe��a��F���� 7@���O�M5��Ń7Eg��e�jS���㖥�hXò$���]iVJp|,jl'ߦ���g��뱬�����~��bp�c�C��/O3w������}\�@��~��J	%.9����}?Ew���hR΃��}�P��#��E�h5�H�D02��:]��9��Dя���~l`M:��i���	i��ġ%��4������a�(�.i�u��ܪ�jF��0FU��s0wI�㶲?� \*�����g�4i�Va�1d�*dVbh�ʗ@Aә8��՗Կy�4�[�����w���7�M�_��zUB���~��-\�K{���߼�s|�������c9��A���9���[�7.`e��4p��[�#._o?LQ��丅`�_�Og��H�V%�o�!"�Bo�V�z��ג#�yw[7���_<�[d���A;zHh�<�H3x��f��C����H�z��Gq�@)T�̼��?8�]3'c%��a}��6��Е&��X�.g���K��(Y3����M�U��ڤ�S(���0���%x+���s����H�f�?gْ��G���+��
~ �6�Ȑ�]�U�r_Mw��r�]3�4�{Ӌ�����m�x��{�|��޶��U>p��b���dx��
Zr�~��Rc�?@y=���&�E�l�U�v��6A�5�ŭ��OF�W���)��S��«��˭�p��EG�OX� T�-�Т͡���{�������MJ�c�yF���5�6G/��ّD��-�ܯ��Y�O��'�z�����ec�x�i�!�>֍�I�0���,>G��7�y��gqK͝�s"�f�y�"��QB��%�������Wr05��P�d�*�����]V>��۴�RCY)�ʤK=�F�[��ד�`Sgȥe�Us��Q�r�I#+�kF;�>��i�o�)FhIǤ �
>a�y�_ypp{�v_��4�U�Z5�F�ײȋ*���f�	kI�3g"�k���������ܓ��Kּ�)9�!ćC!��1��pƣR��+�WD��9��G̗�H��87>�4���PV����,�_�>�x����q�!.Cع,���=�ּƴ�z�#��)�%���/�M�nުis��e�(w���/�R.TƤ��e �`Ԇ*m���x@{�pX����Œ���e��o:}C����	|E����q���m�ƴTN�j����OQ ] �;�ڳ%|8��+_��qM�EH�3����_gԹ�:j����2s����󻂰U�:hfM`dPa�#�i�7�-����ᦍ��Zs/ ��&�'��ߙ�H��]�To�vIY��g�O�q�E7^s�-�ƺ�u�1���˹�x-��@:LJ<����M�Ή��2��Uʣܻ�vX@;2�n�a�G�������7�L�,���ɷ��Ź���Zm���]�yb�8���x�M���km�2���n��:������Fa	C�Y���{�dN�	
�c[9��E�ҏ�n^q�'�8�$BKo{��͂*4E����c�:�%�v��%BH�C �r{���6�!���.�T��[��V9~'�1�p�S�9�&� ⽦A����g7�YI�܎�X��G9����J�ֿr� ��N%���&�{�S�P���B�Ļ��3�"��-�	G�+��}��;��ϫ��
��1�?��!�ȁ���0�
��q�}|]���fH������&>z���ʌ�ϯ+��h�ٍ�*lLE����'�!`�����J�w���b_�h�sҭ����vg�ey��̮hU4�TIo���"J�r������h�a'��e�Fx�' t�E���T�I|�:�W�}�"jP4v�$�!7QW�����t�Vd���cϢ�	-��Х  G�`�����֯��qy-�;Sf�Tk=�JGP٨L 类��ә��בy�e&͆�FB��q���(��δ��a�P<~OE�bb槀��/S}�]�yr��p���]Q]W{�̳�o���(�;$�觓R�q>|Ti�]���c^����P�I�t���柈���VT�舐��f�#���#Up���49EJ�h��A��59S�F����$� ����5��k�1�I��A�
/c��6'���*��!P�cXwJ;�YSP �c�h���WTt�x�-4S��se"�U^���)6�+�`cݯŔ*%�����k�C.�Y!�_!9��;��ŉ�ʃ��Þm��"�O�I1X���EZ�@�&/J��)�  �K��1>��q�6���� [��j;\������8���k�Ӷ�D��ֳaS��jȇ���w�?\oӑi'�%�	e���c{��H��e����ӏ\	6h�  DX'�� ��*2�ޱu�`g�d(��/�)z�k_��$��l�hzM�`��\G�Hf���i�y t�P�hOJ�MEy=��+��H�W`
|�R_���l�(���~3���M��`��\�X�˳y���[��@.��<���R��Z�O��߻ס4r��t2LUV�>�[
�l獓�/�F���'
�9<Fm8������u4�%�nP8�T34x��Ej��^3y��ٛq��n��*7wBY�fv���̯�%�����$���h�q���<��e�\&�sZ�𸖶-�EP�xc�B ���b�<n�7T�{��eYh�Q�gs���FR�(��<1���D�}' i��~��(,x�g�g�c���p=s��ߔW�2S�n;�up	;�`sY���A%�cƜ���,S�~�1E�A)���KOڨ -��@��	#�Y��_w��A�\Ԭy�Pd�1?�'Q����ob3�\
j�F��M����0w.K׶7�z=��������++�Y	*��#�o���q����b��V�D�v7y��Z9���m:(7A�pLu�8d�r�%��(U��B�]���ǒk�Z�g#]ܔ��������9��v7���ٗ��L���K_�j�?��"Ws����!�˄d� L���mM�e��~y9gU�% ��'9��/CÍ�2���]0Wpw9l��PۖG�C��'���n��R�b͑�>w�/�
I甹��뗵\L�=����V��%��F��[^?�y�����Ξ��}?(p����Ӏ�5U*$H�}~Di]E�X֑*"��ġ�jT~��:��i�l�a����{�@�t4<�ߕ���Z��Y�u���7.�j���K�U�6s0������ W�UXG�";ziKKa_�~IV�GNe^A�3��/Y/���Ty��i4{r���wꧾ��PM����
�B{n
~ aO-׉ KVp����c�X��C0�N�/c�A>�9[�[�g.�ef�<*��V�~��o��$Q�<�3��`�oUO@r��e�%�{��|�0��V��e/##�4�[r#R�w=�V���MÂ;�5�/�P�Z�3S]��$��G��}L+�ՇG,�))o߼;ĕ8�nE'�Q؅�0l�1�,�+�;�*�.�� ݎw���3(/�蟊�⥳�T��8��K�%�n���ޮ� ���aW|g4�f/��ǈ�K�vۙG��]J��m�w����O�p��g�f���/�maأ�v��|c�h뙴e�p��.�������m�rxI��M��?�V����0�`��lc9���b�q��5FI8���{O��n���!�#$N�f���щw��E�~�XdeTz		ËA�����K߻�vB��OfJQo'yAb�
V���p��:=D�������]dw�y����'hzzT�h� �ye�ƞ�DN�ypek+�0��,���w7y��q���N�fJ"2#�Q=�j�C���r#!���+e�e���Y]Q��6�R��/��=^��[�� �O�l��u~b>"�-as��kQksI�&k!��>6s��h)A�m��|��vva���ڿrpV��_����5�RP�T�*��3f�צ��f3B��k-��͔�P��D��7�K�>�)T�S!~�C�[3l�s���M?����0W���9�J���uH��!7y�@�9"��y���+j�z>���u	���AC���5EI���F�%�#�����!�e��E�
Ū�]�`��w$�/i YI��R� �x��Gm����|ҏ����+�R�ٛ���_(	�h}���>H�d4G��������U�������}h�_o�|H@O����m��١|�!��x�笁�E�b;���_�➲�CP���O���1��H����3U��%haG�d�V���4��R|0�M`z˼@�=�Z�	���&'K��TΉ��D=T���Qc�RֿDLD�l.7����ǧQ���}uUG������-H��@5�.<�����5���z�M�	��+�v���2Aaa�mn���ŷ֊��g��,B���Ҝ� 0���+m�����b�T|���M��kH~����
	l���Q��:Na$��YU?�{���N��
8w�9 g&נ�|�`�Uq,X��fÀ�]'o�&����E|&�羡�:��=vV�%�C�®{|��Ѩj��˔�m%[t,�9�fG1e�nSū�&W-��X��<o��W�g��I�0��	YBXb��GtR���L19����m�KN,:��|���C�S굢C����C� �3��.�	}J#+�E��	���e�����?�6�!γ)�y650�(�:K}^P��z���{��^�&YP�Ddj�x�@+<��{�Ǡ�l���*| ��隯@����;*�:�F��M���_�Q�.�4��xK��@�y���U�uP�O��o�C�X��0��KF�CY�b��e\�Sx�g�t����Q-��'����A��&����6j�K��z7��^��Pqяdq�຃&���-1+����G*��ZĐ��r���ԓ��ۏ:�=E8P�I�L{�3������@ˑ��m�@���>-&B,��q{'���ǉ��|(�<�@��=�Ч����}�IY+�rd�����]̙�{�~K�Ŷ�6;&(��$*�s�qY��i,���s6�^�u��I�A��a);�C�ځqC���ǐ�.��a�j�Uk7���ЁJv됆\}�5�1:S�
���.�� �"e��� kw?�I���Als�c��)6b+0�ź,!K��HQVw�ZYn /� �h[^W����n-/L���}�"�@^�u��4�+�trcIf��/���J��'�2C�m!����A;�6� ����-֗7�%O�1s�����a@��/�1Y��	�e�˂��6�60��:��9k;���8��3����c#��_;���<�b�}��U��:�o.�3'� �	���h���)w�eAe}����J*dP���elsD���۬�"�uI�ˈ_�m�j��j��s��[0��穾S�z�O/��U�G-�R�z8����toX�Cu]߈&�=>����d�W���f~��JB���p��O�J�TMb4b`��}\.�nש�$B�����^�	��RY�ʁJ� 4ѝ�\Q���(VL�G���d��K����/c+�G�l�T��m�N�����ðAf%�#�8Ϝ�4�Y�� ����9y#X��LVn��*ҖfY�y�Baw�F㝑���$��'���������Pez��� �Z�9�э�E�P�c�Λ)�������x{��`Y�VQ��fs�>�F��S(1z��Y��8�i��W"�xt�gʧ�ŰL=n<���uY2�<]nV���M`;��s����K��^��X�kS<��1`y),�K*Y�[��ە{	ZӧxI�_2�A8���'T�P?�n?��3���.jD�f�=
%q�F����L�K']��{��`Ǽ'��+���	E����5#��m�0� �l��Ɍ���l74_Au���(�(l���uz�1�m����H��~n
xaO�B� �5m�#�m��V�̘`;�����-T�1�c�l�'�v����}�9W�1�>�z�M��8� �wc�S~�Mk�0�yۉgl�>������C�z��h�f�%Yw]�)�prf6l�W��Q\*�&����0,Ӳ�+��b�1X�9oC/;�O����\�2�ϷlǑ��%d�����?��ؒJ$�ι��}��[���cӻ�5�dH��DĪ����#:��:؟�E�~��z:O��i�N�D�A�i|��[� 4�i��Ð��C��dj�u�(�ѣj��f�KU��s�k�YIP R�'���ԃi(�a��Ń��V�F� E4A��ߊRi����y�Z��ǈ�3�w%�a�m�!M�I��0/B6N~	-RK1J{�����u�͓��0�c�NzA5�M9�0B[��.օ�c�����To��QZ_䮦`��O{�d�~��%�a���L����V�*���_#��[�Yw�;��Q�8̨�D;��J��2 3.�{�Q��y�n�x�)�0��G�B�)�K���8��'ٝ���~�,�x����A�.�Ǹ�	Ķ���3cfq����ݷ褯��k���f��43�}��BX�B�W�\45g�ke!7M��m�Ư���h�>Kg]�^��h�`w=(���8Fjv�qLx�A�!��m�W�q`�|��(�T�ɋȣ��3W�T����vr4L�H��?�S9�b,��{d�l��^�Ȼ5׬=�5ឣ���QO��mޝ�>�P��O��g���8E}?�X8�T�\��F �����q�/�^����2J욈y<�e�*Ϭ��� �0D�D����"C].��X4'�#9z�2�j~eY�0�-ѻ�*1-�0�֪,����@�{y�j�qA"ȓ)FfC��"͏�Q8���ۄD��y��ex& Z�H���Q#�J1]L�7���R�$z� ߵ=��V[�n����!����]�z��sB�AQ*�	IBtk�0v>qY���3)<
��Z��X3a"��U&�p1�_&�$���B5�~��h��*k�1f��ga�E3Ākh���/z�����IvKL�)o�B!���C��<��Ҧ��Hٟ�ՂW��9��̍�EHd�7��@��{�PǯG�*%�_>�L�����eCN�X��	��Lc��	�#^B*�9���ʽ�����2ટ���[ywp�$/$��d>��� ��J͸m%"\�w��.{����P�Ieň���:�<�
}y�ݐ��r����w���O��cj�0�*�����w̥O��AD� F|+��᰻���E~>{��g_D��=�����(�!��,��1!�U*�hh\a\d��ә���m�����H˗��x@Z�r�����'��B�����K$Te͂�,�ӿ�K,�h?�g�f7W���B��u�|��x�p�/k�-�|�@0"�<U�������҂���6���5v�6�2�3 aǳ��L�뷑;���YB,��b���;��G9�m���'b\����"M��_k#dޣ5B��4���6���a?_YР�{�f�N,B�
Ӫ�9����x��qG���ڙ�o��+͸G1Ew���S�:>��v"ʯ%8�C֩�{C>j�l�+��w�
JO[/�9��Y1���S�=�&�����o�7w��	�g���I{�܄�X=� G�*!�1,��(9�(g�NGo���`��+TSY��=���^s�q]�3q�1N�	�m�+����������z��q"H?Gʆ!�ٴ���0�f�uD�}�~���� �?/�� k&tF�տt�S��+w�`��k���l�-�鵐����G�u��MD�����_8[����D�l����BîU;��Jfo^͢������������C�� De��=x���tW��x\�B%u�?'T��R��!j��Z���7L�&}Ѫ��d�B���Ä�?-��ӥ���G����%���ꃅgP��:�ʀ�=�E�P�
�Lև5�f�˙ףƑoxճ2��y~�B�p�qv��ތ��D�۩�v�<tRI��j��O�e�;}����a#r�d�*��]G��{�j�� "щ�(�̥$]�V���qt�6i��E�N�p^�_�FI�. 缵�������RS����p�܍����Uf����J1���ww5/o�S� Y�>p���#� ����`k2mVI��A���c�$6���`�a!Fj}��^�w��zY��E���h6aiWʐz��UV-*e[�)�A"K�M^�0�S�+�bc���ʫ��
.aԂ~C�k%!Ƌ\/^(;�ϭ;�<ʹ<����z��`O�k�1����;�k@�-�/��_�i��ڧp���lm6)��:��(�;ғR�ӹ�.�ʬ!�!�?�z���~Kjg-��R��Ґ�5�o��'\�		�Ü�n�tn?�Ee����%����Җ�������ۇ�c(�u���Z�ل�9�{��7����[9�i�޾�؃z����ƜG�I��5����t��l�� ��'�=��+����WaM�Ȍ���H��qe��@�녫M���`�М\w.�)�ө�ա6'��ĹO�D�R􆒁En���_�������LK���ѫ���.���덉��/u����Ӿo�=m.�Ջ����n%��8�l4.�㣻�@�ɒ�y�E5�'�WnS!*m�BY٬����a��ڑ�$4���p���p�r�eu�r��DZD����aEF�gc��Yw��F����{U��Y��^QOqs��F�w��+1u�ϴp���iO���;�xO�Dg��K8�=i�1�J��2�F�nq;�f��;êVs�\f�w���Y���h�S���1{2)��XK�����vW�	Oɧ��|_��RAS�*ԢN[PF�?+*�,�e�����
��F�����#��@�KM����L���ż��z+��	`}=�'#����k�����������7�Z���z�(�Y�9u���h��@���9���$�ͽ���c�#�J���	LєY��S�L:?ٍ�`�;��I����P޹xm�W)���&��Ա�Z�� ����E�M��t]6gǷ{�����/���]�C���`+]:C�pm��l8D����Aֱ��Ӎ�Z�/�bA���4�r/`M�
�*�!,�\B��ت!�̢&%�����T?V�M������}5��~���th5���Hٹ�D���$��>j���� .E~��:ꁶi��k�rn�$ w�v��42�C����M����u�T��$jw;����
U}�Is������
 M�5싘�QiCaU郻��Vf��K�A�����k��FB+y�6*�����w`����M���srB��~6�J-;�KDK�:��D�+��w��Ncj�AP��9�%�[^�/.���S�����4�.op�<Q8�I�)�]`��O��4��[%�g�2�sa	V�,%�#_
5[���X��Lw����;D<eaG��m3	���
�9X�sdD���ZG���)��{�1��8��y'
��2���'X�����-<.��݄0����O3�݇�=����y�
H�&R\�Bp�d��$��$ţ�݌�W1jg�:�^��ڔA����y��]S���cW�w���ʎ����@��5��r\@�m���l��|�(�ɦ�i�$���v�ζ:��r�>�Cz?QqG��oٖD�lY���y���5|���#OW^�(2��Y�[�\�e��!pbE *X,CT0П��~��j����9���X��J��!y7�C�rE�g$.�]lDy	���[e�]���;����'�Mzʙ�6��e��.��+�����N�0�+�,O���V�y��q�|/���f~Ʌ"h6Q3���6�>���M���w��E�����A���(�]G���3�Rt��,=T��[un��Ŗ*�1�X��v��s�|QE��I�}�k��b>�_��Px�)7��ǵ���sa=c�Ь�pj_a���&��5��r���E*&,�f�P�]P3���k�����j���ܤ�K�{)��y!t��C�����A�wC�N�<��Wu8�9����W�H?[�7��4�o�W����I*��H>��P�kNF�ǙC��k�(����ۀ�#����~�[ȗ�
�{/�:�VR�w�H�/߻�㣤H\� z�� ~m����r΁��H5ڡb����"��Ew*!}%���Й���2��+���KB��7��e0Y�;`v�rp'Ob*�Qо�+�|�T8��	:�"J`E:��֔_x_��kW���g읣p^��0��l��U�YhW�dda)��T^����n�C���rSu����ZDD����'4�����r�T���������z�ҕb�a7o&�=�
��auK��S��j�-~$@+�+<����~DЉ�b�C��mkv	�2UFwa�E���q�L왝A�,8~��Zh+�v|}�ⶶm���n5?b��� �OM��&k�i��pT?N��������aZ|YK":{p�Ng�
n��9����V��c�qb��߼���Oo,�3�S4Er*��t$N:���v=^�%�.�C���{~ ��d��e��eFy[��9�D�1[8�S{�&����?2��1"gh��I/�q����X7�G�"y��+'�F������Nb�^�rYl31S������J�����Y3,=zL�K	s��+��g�:.�����u����4?~!ꑴo3�0��!�]?}M����������^�&�\��:���.�r+�)���=�ʊ��;v���БJ�%���5ְ���Z���B_��$�p���0W��U�5T�}��U�XI�Eͮo�!��a�þ~�
�;��L9�E�e���x�G�t�c������]���,y��o�.r�j!�`�Ha7b��M���Q�dg�	�p#3�S�|-g�����G��>�Х�� �O���$��L��={s�P��bL1���!����&ʑ�^I����Bb	�qq>\9�m��_���<���$��1�> ��}��r���EA�]�r{�v��;�"l��(��$�~���$q��Ci"T��)��^B��}>I�;��b䟹��������~�+ݠ9�Ua���E_[J�P����5�̴S�؋y�d� �H �F� k��I4�WAb��cd�X6�qI���n!A�-���rw{e�Y��D�ޱh��WOb�I�5-%�+τ"�^���j+upFc��N�e���2��ݕiC_Z�!�Q6��:;��v��T����[���ZOE��1�9EĶw�@���/�Ͼ��z"�3���]��' 6DH��Y�h7�;~��n땰)b(�|�+�"���)X����� �Hᢵn�0No�''Z	���^$�O�7�Ee����� ���Q���޲�����b��c��uX�Uq|�#��Z��R�}�Q�t�D=����z봩�W7G������e��9�t|��� 4��H�=tе��Wq<&�����g��R��eQ����^M�{�`���\���䎔����S�ßu�2R����@`�����~����L�iȬ��q�=>���_$/��)��~>��ym����p�Y�&��%��8Ō�4�H;�vb���\?ySe�b�n=��*6�Y����������[�BM$��ʠg@�"V`���ep��7�=Z�*ʖ�E�w�c�z������Cn	�H|{��Y�L�Q�=�sm�	F��4G1p��H�����i9ŧ�Muux*Bg@�h��C=d�ߥ$2Ip{n����6�;���s
�����TD+��S�<�1�~)�IK��ћ��9o	d;�.�1_�1�An��iuP��?f�4��OU`�9���
��Fݣ���UK�gD�KK�����ݎ�+\s�	{�y�3�#[O��C�����XdUy7� ���0���(�!��c^u����c������%���8���x#�����Z�X���{��y�gC�o����%΄���;��sDW�~O��y��j(���
 �/\��,�M�q6�o�>g"���Vƀ�J���pF�������]�|Nph �l�PN��k��\�4��� �hT��j�b�Z��/�=/�P�����<��\�v؅q���%��7��i?�@��_@��zC}�ᗛY��1�5&:�Hԇ�Dz����]��Y�N�0_`����~Xy:�g�i�`��*��㺡��4����po�MvD���\u��4HxEj2�ɦ���U�os�M���*m� H&�i|�Sh�i^�a�CX��i�VN��6r�A��{�@�}��ly�2{����c�w�&�գ��Mó!����B���~Q�-H��K�]+�ut��߮y�Ó��_/c%$�AkTg9x;�[9V�.L&����y���WIo+��QS���Gh`^_hO�SY��}%��Ǎ�b.�V[l���#:%�[#&�H�\�Gh��^�H;�(@���(��3�N]R4�¯�Y�n {���hG]p�)�'��(�8aa�'O���J�"�ş<o��_>.�y�����W3�tr���:��;g�e�E���1��Þ����_g�xvG�RNgE���!5%Д�ԩl�����2]���^?�w����I�u��$�g����	��wm2���g��|t�h��m`�������,�Q�6�uW�rIif�>�?�����ݥٱD�l���~�,�"��5�b��F�O�ƴ��"�t�n��<$�b�5�\I E� �X@�T�c[üݬ��@ҙg�T�qe����J"R�y2�B1 �"�`�6�D������ݯ��|HꟅ��'y�Bz��r�Q��eO����JA�*��<��0��e,�����y#y�q7�"�߉�f��A"�rQ.���X�t����I�ݘ���R-�@a]B���G��R/pێ6�@=��8[P�ۓ ���̝�S`�э�s�PQ`�I��k���>煉��e�)2,��^��y8aX_��KS�p��_��d��D�5�6.��n*�f#bWO�3���k����e�J�|���K�)���!��GC�_�Z�����>� ��8�W0��9��ṽ�*H�}7*�
�J�֯��)�~5>u��� P^��C�nե����\p�6s#�'��ͩ���pLT�Z㲪�q�Q��w&z/�����(��� U�b���m[��m�ć�5��\�y���~զ��0���}�j���ɼ�uM�����F��@��ZƠ�/���m4�O�m���F|�����h�]�]E�U���eH_��β&�}��&�绋TQ�?�U`��hR��d����#���0����*�M"���t�Z�5�����'\��߅]e����T[���p���A��]��7������&��u�G��.��˥��-�1@&xD<�ʫ9��������H;vD��2�x�a��z�CX�����It,��Ҩ5���R\�}Tpm�=�ɥ�b�g��;��Mv5�kُʣ��V�%��&bM��kJau�Y���{K��N���
	r9��ױ������q}S��+��q�og����Emܥ���:��vXe%.f�C��{�"�ݢ%�����b�[���9��1ֺ-SV�^&��)��-睯hx�g#߭IJo��za&X��G%;�gK6:�����N}9���qG[^S�d�s�a���f�'x=3��g�	�D+i^@�u4!�R�>�p� �'��?�Q!5R���m0^B!�.}����v)����ꏽ�&���յ��	�+�mčL�ˠ����%�1����;�j��W���P3�������_��_�"��<��b��Ѵ���W�Uq���@�so�aai�޵���z��v��
e-��x���t��m��x�6�5RJۦD�i�j�R���7��N�2a��d���K�1ώK-s7��,`G;vߚ�F��;�]�O��>��@m�=�WP��$L������ә�Ցeeɳѽo��<B���ql
!��Ǻφ��r�<j���Υ��lh��!@}��~j.�r�i�`��]=}{����vL��Z(�p�$���>y q�L�i�;�[>^}��Fw�I�hb�r.9�tV����=��̐YTbR��;�XU\����V�J�3؆���5%JtSe:�������> ������k�(�IO��A�lAc?��6E��
T!<f��Yِw6^�Y��+��zh�F�W@-���- ���߆p"�kV^�`+P�c��V� ��� V��89�Ci�!�78%�y;�a%�����q���x�H�O 1�
��1lc@��/6ϯ��a3��٧&W���D�6_����Cf;H���	=��$����5������|�t@Q����V]'�P+
�+�4o?R'�P�	����)*X`4fPeN��ݿ;�u_��W~�[@��0�=*����u��PW��~d]����mKX������%pz��k���G>���kl��st�2��Ԧ��9��=}���xVW�7��>:[�0���Tӳ@����#�M3O�`�>�\-2n˟��2@ӡ,�u�zQ�����R*�*�;rlEe�׍gK�2LA�Gȇ�4�GӬ��Ѝ<(/+x��x����xUm$��K��a)�%T@8�44�ﲣ1����F>y��A��>�nx#(*��#Y�r�Sx��w� �'�$N�B��]٣��ek����Z��B�"n�E<;c^Nx��s��|���,�5�{��iY��1QL�sHx�F>�2$�z1k���j��ib�iT[���ΐxˡg{4�ŁoP=_��� �)2�0n�?\�;y�sE�eխ���O���i�jSm�1��)|��K���V;ڬ:�	�)��f�_c��A�iԘ�P�9�?�|S�b�L[��w�l
V��F4f����zK�7���F��a��8��+�	��}�o#6/���Ĳ=?���q�7e���1�pB(��|�I�uK/j�^r��i�⯱��
bͳl��Ʈ#I�O�'�Ř��Q�'y����nك ����ο|���7]�n;�W�T�oJ�
D��PΟ ~���4�M<`��j��g}�����exӥ�'������/<]p�;pc��l�|�ۂ#�w?����C6覥�bw<�*�/���A�W@�\8T�`��B�>%5碝~':?���{-��
 �}+
�4�r�l�5��H�u�D�RS�D���t*����"����~�W�: mhi�[UH��ǂ��fU4(EװK����}�5\�u�<��{j�����9UsyswSF�
KI( Cu�@̋b9iyO�aK��qM V��Ѹ�A��rߛ�W��+�y	OQ 9P�>�Nw֐�>W�M��$�A\1Bg�1~l�f-�s#K�����z�_��C.����cྎA�F�9�p3[;.��WꉚC�����1�o��dQn�w��>`9�O,�ѭOp�%�ӿ���3颈V)#���#`9[^������By̹Ċ;�d���^��m3�4���A�J�s�i�͏A5G78)�Ÿ�'��8<�n'�B2�h?��Ɵ���r�.���zi��oD.3,1�TZШέ�������S�
[�Z��r�Gޚ)����M�Hg���R�P�M�7�G!-��R�]�\
�YG�wN���C����┴������&m͖z�by�|��������N�]I�,�:�r䳷�99�?����?��d�lOX�YP�]�75�_�����OO̢�9+ޏ���R���=�?�BrENA4X�s�T���w�~�	7��q)��YюΠ�J���y-�}v���WW�Q��Do��tc&������\��V3'��z@��ln�e�Do����eM��i0�5},�q�ay>0"q�����snf��"��GQ)R��B��/�5���n�p!���F�Q� �x�]=�#��(R�E�Q&2=J�[[+�d�;�8�g@�NV�,COss�Q{�<I�Tk���>"����sd)-���k>_�e�as�'���p�u�_�6c�\�S5���y�7*��f>P��`�3�&�kV�� �c�n��ZQ�K}��)��!jR�ChK:X�X�wh9O��W�1'9����?H�h'7e����H�����XB)V�&>3���a�9+2C�뱥�i��a���z#�ʹ�|�Q#PK9��kj�p��L8tw��/U�\��u�>M� 0}�&m��3�hJ�?C����0Z2���b��sA�F�}J�l���ی�UO���aً�A_A�5����b��q�ݱhO���M��a�#|�o�rG瘒EO����8_.\�����4j������f������U��ChMo�d|���c���M�9�=�(k�)?�ZzGቌ?�'��`�@Ͷ�!
T�L#н
��>k��~��X�+7%%���T�AL�uAݔ�	1���:-��	@!S<f�:��/{�#�j�9x �#+�v��2���a�E��]�������q�,.��~z��H��"mܮ�$6�b���V��M��k�՘����uN$�%��߃&)�a���YA��{&ٷN��
��9��e�̧�L��q�<����k�o�ÿ͉�AEh���*'H:o"vs�[%���Cg�{�D�=�?�����[`�f9��1Q]0S1��&C"A�č\(Oӯ���g�1�Ie���NuX�PG`sť���D�9��Y��N���h��"��S
a��.P���*Ă5�3���n�	i�|+DQ����������k�t��{�?xE�!:��e�C09�&�}��y��
�P	c�J<�&���0
����d+(�>����(���c���-��t��M_K��&���n���0_I7�z:�i�ݔE�S���ѾU�"�;��oo*��D�����"� ua˯�N0�e��x���th�=��������ہ94��r�jWꕙ>87����g9���d]���&C��ɰm-�u��炖G����F��6��؂f�����{=�.P��L��;����(����U�����*2lB���qg��n��u�R�� !<�F��FZ��$�6e}�e��CrPf��{S�]��D{]�g����5(��w$nom��e q�ЖiC���Q�^��ᐖI˵M����/΋��?uD<�4������"�UW� ��m�Jb68��%65���S@�f���q횒$ ����� kc�Ij.AXU�c��6N8��1e!7#��Fw�v2Y� ��%0h��+W{+��F�-p��:H"|!^":�nc++�Zc5��ś�����Vԓ� C՗%!>b�Z�;]Z���ʊ����ї���O�8�1���Ĭ�Q@b�x/q�t�0h���c��pV����6z�!��B�+;��ܝ����W�23@O�+�˗)������摒�����&�o�~�'��f	�ȵ�T�C��o��e��ݺv������<������:�z�1u��͈K]V��)��m#ш��G�����?{�zT���`G���fg��  ^t	��LK�t�=�a���W'S������K���uL��d�6�9M�B�`�b\�x��Z�b�M�>��J�UM�� �R�B��6�H����H��9�L�e��b@ַ�U�s�w�z9�/�)�3� ���-m��ŋ&XÜ��%�5�8���4?�J�짆�Q�y�ɛ�;}n���*>U(Y���j��2*�B�$|���pH��|;�C�4ef}��OZu��=N
E�9c9��
"����I�}�{�FuY�§Qz�s#v�FyC����1f�����$Aio��CH�x�s�g������=Zx��[/�2�#�n¾�ן�;TF`s�j��Hf��J8���d*S(\1�vf30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�/ڜ4�{^�{]�$Ht�E/Z}1TWZ�i�ˀ���9��Z6$�x���<�������5~��ߣ�L�8�6Z�^��3�B��˞� �Z�>~� Bc�wz�荏�`�ر1�y������P��v���cz���Q�ا���@�j�{��T�,2)��2{#��X�jEǁwNրv�t-+ ���2���)D���?&Ìw��K �ڀ�-���9E���YW�%����e�1�8�3��c��<G��Y>i���9+��=��in3�4�S�@���`�����j�@��I�`�39�Ǹbн�>D,:t��N��@wReb�T�
�1�掚l�A{��K��ү�!��'���^g}h�2�+����1�V"5K�AO���9�����sǑ9MܐxZ:"��?�_�=�h���G�9��eХVN�Ѩ��vdv&r���C|�3��|�C�������� �W;9!��&`�6v�8j�����.��kn�	�M�6���V��.r�{h�B���ءz��9�6U����H>��gm�L�U��1��v�Id�}J��y����]�M-��_ߐ�����V�"k\��5�:� �h� l�]Sg"®d/b��..L7���4��GEO)����P}��:�Dÿe{7�-	<~I'�����8h ����~De�~��J։�e�*u���@��2�f��hV1�{�Q�b]r�&���W!��w�/i�{P�WW���h������/�p[��=%>��2ט���i����~���������&R�1�3!Ŝ�`�`�|Iu�i��a�� ���R�>��l�d�l�}d��V����]>��g:�pM0	Eqyjp:��y�<A�Q��d>ۦ��V�ROg��Ayqd���OKwj��ƍcS�l�T(e!L�y���)(�7�D`4^����S-�ة-(�@	�d��-c�!n��f`2�g��<W��Q2)��u����-�2H��F�����f7��J�����oc�j.��	"�k�7uS�57E7�4eY��јIm��<Ǣ�0���ȹ	hئ�����W�n�p���j��&�qO���2����
n�uS�3%�F֑�|sB�K	gi��P����@h�E���̳��h�C�]���10�m�+Z�Pe��5�"+rYM���#ZA5�g��f;Qo�?�3�;"�U�2l%4���+	2|�TI��M|o��1t�PZ��j ��1Iu�7
�8|;��!�-��	������<�7�7\IL��؊�F�oi�#��$E�����`+�ӽx�L0�	���o#�;���ou�4�m�ݞ�>���0�>aU�o��p�u!�Q���k����(��K������N״DCX28����f�j�5�$��;��� �E ��9���w\�)��h ��I�r����b�(�¶6vo��U�7�>�V����P�a����;�U��lTՋ'V��i>� 8#Q�4P�~�oa-�����9 Vv� �l5���2{�����eÚ �P<����V#*�OT�uT�a�ӂ�te��3*�>�7�=�64ϧ?��w���{��"W���B���r�L��m�_?cλD��-���Ъ�@f��%��L�f��F��ހ2Q�W�]n-mB牻^�#%��Ïj��� ���!uq�y�ˋ��5�>���{�� 2���TNO��dxC��E��=`��8�P �Y�%�𛒓1��k8\Z%l�;�M��3{��>��;ڞXs���\(��Z}=��+J�l��>SJ������u*�������1��;08����M�3Bࢳ�vSY;��F!�%���%o���*��o��S�w�ҴDo[�.\�������l �?��h	L3	*�[S�u���*�YjJl��5��v�';h��ˍ�5��ԷY�B(�X��S��5�l�
f��M��ڼ�^.�͔��'���Ԕ�
s��� =E�
��\Ja�\��U���۪
�ayz���&m�� ؍�Rv��j�m���A'.��#�:���c�:ľY�v��[�{�i� <@�P�qM���*_H��<&������D�i��о
�����bv�9����*��d������b�To�
n��wZ����2�*$������<�x��G`�~�5�1��w�|qf���Z���Q�������`�)t��UҞ�]���WC�?6Q���i�#�i���+� �,5s$��P��r̠�&��kz8���2+F���w}@�.<�Kv��F�\�8^kr](4�ʏ߄)稜��As�({����{�d3��et�['X`�oe��>���9Cj����ѡ�l��hu��D1���pLGc�W�z�����ӑ��H~&�%]\NVF#@��n�ƹ\F���n��2t;
���f��|�F�vm+��XT�owE��/�AR~��	tݣ���Eh����mγ��~���mQ��$��2�w��>���9|���m�Z�2��?\F�>J��G����X����_����x���
T�y;uZ�G@LHK�3pz�K>!����)��T���l���g�+����^JJ�!�EfY����}�r�����q>��,�#�����cߏU��̩��q���܀�qM��o7���S���1�\�-�W��p���F4b�F�C5t��q�������즞� ��5�0gH9bf̍�5�?tJ�����'�ݖg毋�޴`����@=:�� ��J	����qa�V�NO/-��
Fw/��7�+!�[m�ڒ��c):�d8��^�`�#�t(��GJ��p���wcz/���{��b,t\%=I�~S,�p�-��mF�|:�ab^���P�˿=Ԣ�_Zq��bc42 �N��#4ʱ�/�j_��{q��$�y�EC���kg�i*{ܨݴ���v�n��$^Ҧ�%{y�:o����~%P߷HY��֭6naÐ�HB���2�ns�~aXc��U�|ԯt>��E3Ky����k�$P�v�NzC�w�(����e�S�;d���H`jU�/�h%�2��0FmX�!��jY��w��v�P���� �2mp����DEd��S�����_�en3G�A�%����Z�Y��`9��u�S1*�̎���<����G��vYҙs� 1�+�{����p3�'_4zL��3�t��i�m��@-�]᷌#3͚��vQ̅��D@P'�~�N��@� ev�Ҟ�r1�;G� �{��������Ifߙ���;� ��h2�(��vo���V���K�ԛ������燖���Y9�{Xxn���x�m�s�%�������͈]e�v�N�y�!�GnC,'����X��� ��+��N��3� �`�?F�����I�_���j u���t@ެx#uɸv��.V�J�G͢0:X"���AQ��O�Lu�:�,4G��FP��O�#� �4ʱg�m� K�hv\��}�F�O��T>Z7�d���^�w)v�B�Ǫ\�!/���>�I͂��'�f�)-�kn՞��ޟz$p?��U�����A>Ȕ����L�[�����K��$$U��n!���~�=	���5?Ԣ����j���K�X�ݩ�R��֧�X�h������Z8?j?��/Љ|����a?�9��TA�
᜼d_1	Xr#H������R8I��[��i�/ V Q�5�I��K9=ȑ�[���(_c.j
�`��k�6Tl�j��6|�m�0�J/O~y�x��3��k�.���]C�[<u|9��E�I���Mx�4�K��
D�i���j>$��h�E��l
��`#G�c�'����,Һ��7n�zWX�=�,)��M1+0ta$�szq����%����º�+,3�ћ�;q_D�"F�>����.��G�k>Jj����'J����o'��@kV%R��\�ؚq�*{�i��ӲB�X�2%w�W���ɭ9���QD��E��W�r$wz�0?:nY��n�4�vr�K�aq~-q��W�W:��z�p��L��P�OL攈���}�M�M�6�8َ^r�4aŊ"���z��9�^~&3_�����O�#a}�ʦ,3���)G�;�R<�~��i�f� �;��HB�mC;D(��΍ōn=L�a?�WV�OH��wm��oڝ�39�3'�����jf"A_�g�?�5���:�y(ip������9� ���SҔ��WU�:]%�{��wK�A��Ӏ������U�'��1���t[]�d��m\�"V%#S����"���ޛ�)w�5ң��+��V�>;��h*����Ӏ��uqQ⋨�E�(�č����"�}��a�&]��y:���B�A���F�
�Gd�H��}��Br�dO?�NF��WK��ؘ�
��doq������Ĕ�d�S.�f#WPQ\^Nj��@z�%81���\{dYS	�U����*�
��>��18wQvA�x�IV��W�>t�X�<�ã��9�':�+�����w���Ȑ�;�]i�k�V\�\�&�Lq�Z�=�����	\	lr[�S	7�L�E�����Z������_@bZr������#'�\�F�����y��Ĵ����P1�噖�pZL����c�q?^G�=i�&��3����V�skK���M@s7 t[+&03�8� 8���W�*�(��!�ps�������D���CjuM�����S�FBҥ��6qRn�۫�9�M����0
r�Z'>Ӂ���ڳ�?2�����>��:�4f��U*�'��,{��y<p�1�������4���f�ƘL���G]8�cL�=FQ��:��R���۠�jܞlƎ�w�sǦ�r�E�,qu�����߹9��l�`(g"-�r5���Y���b�-�����gz��ٸ^B��#�x��7�z1�O�����'��_D|4-B�Jާ��Tk_f�;!���n����؏s��3@�?� ��i!g�*1���o%~Af0;.�cg6���2��Wt|i�*�(�z;�
��G28Cz�D�-��fY�H�E�r�''�LPG���P�C��I�\{�K�T$���
^(TP5�u�$���{A��n�����sU-��4P����)2���Mx���Zw
��Q�p�O[�>��B�%x����D��W4<I�刈�p��_���\W%�:>���+�u�}�^�\Ͽ<K���)X��U�i��"bګ����>�^�x�C��p}p���T����Y�	��ܷ70u'�vEϼ��-����b5f��XX�n�[J����m��N��j�����J6NW[o�V,/�_�:�� �CV1�w��$�
�4�ldܜ���@_��dnD���j���?9l ��jZl�<�/3��E_��ѽ�Y0N'u�93�~�A7���0�}��> �]u3�~�تg��k13 &�o�̆h~פ�C$8e�$�	��h
.%�_ 䕆Ek�Q�/�M��{zI��[[��߽۲��K�Rٌ�؝�c /H�iz�0��+��rc+��G�C����U��+5�����X����9bP���u8y3��f�P�E1E9.�8��B��;���sX�
��[�{���|X�	.��n�<E@H��_�Շ���X)Qgw{�ȏ �7��Nn�=�U*�@�W�c�c���a�)�/y����<�3û=�UMlF�R'��\&e�m/Ew��ͼ���6G<�� �ꓥ$�<���]�.y/���4����;��@$	w��:��<��_�W<Mί�x��@�3�5�	#�N��X�wB;Z�e�?G������{��ӨU��p����5ӑEKB�+�h0�5�V��%�x��n��iT�R ��������H+J��b+�K��*4������)��?L��J��(��I?\���`:�R�\ŉ��ۘ�QO��a�(drYq$�]2��"�T0�I�	6ѻ^
��[|�_�d�q�s��E�C-�U�DKI4�LU��܌�� �e�/��@X<�5����K���N�ŝ��G\~�%�Gcf��X���} ���k�IO��s��̤P%x�������^�]��W�I�:�����q���}c���x�-������(��Q����tϞ�A�N�_�3llر�Vޞb[o}��f�E�Ƕ_٨͢�����V*B����b��Nf��<K���x��d�5�j�#��a~�v�c�u8ݭ&����F`��Z��Ύ�F��@M弭�R��i������|�D�5�R��_��|^^�g�D�2���)��a,��f�L}�t!MT�2N�g���ln\E������A���Pt��}e6dl��J�"��R/��AѬ��Q?v�8\�r�%��n> �Ki ����?��({����Ku5;J����m� �,���`�6���(�x�M���n�>�ӎ�jo?c��5�bd��MǷ,�����*��PgC҂j'F�q���73���0�q�.��'���$�!4`勄��.�jDez���I;nՎqM�=6N!������{; {U���j������v6~aHH�g���Bo1w}Z�v��Jo���~��'0�]U[8��"L�p����!s"�x��`�ꍆ��-�}] �_"oR/Owf.�5�7<踥S��u?hO6�h�[@�A��D�&�e�Y{7!<K�J��m�E+�:���^^uDR�L�(�ֶbĵ��ƞ)sn�?5EYTV~<���b�|�ζ��픞�^�<D�(�Ϥ|�y�ә��P�'��p(�b=��|�?ч�zX�kd��Y����1!����R!�73.|7�yR�����V��������� T�R��v��KdQ
��(Ŭ�k@�w<V��BI���i�q3n0v�y_�:�ì)�bQb��>��v]�u2g��myU����Kd���S��S+�T���~��ܲ-�4�7��f`!J0�BSI���v.=��#�d�mC-M�n�Ky`B΅��:k1Q��Ժ$�?���=-������ͬ��������r��ܷw(̶E�k��n�5�2
d|��YEOP�V��d����Ƨq̹��G�ɞ�dLPn0�/� B8�S�k&�䳓�*2pL��� ���s!n\d{S�L������(�8��i4gۻ��s@5��9�B���	��֪c��P����'Z��㹥��"����*�x�Z��*g��HfȢ�o"�� �p"8X��?�74�j��x�|�� ���!o��t^����� ��I"um
Nv$|(��!;���F3����[y'7�I��*�%y3�`��q�#��q$.��og��m�K�&��0�Q2Ѩ�#�2M�c��u4~/4)���d>�R�0�#yUW�c!��܊{IHk��Y���>��8�����[X��fp�w�u���;k��\����f��D��)<ߓh'���O&r(M��Oi��O��v� {U�U>�@̟��\�����B.��(�TP�ȷ*>�'�#^�JP~ao������9�	j�M��Y�ݟ��h`ep�C�_���m\��#G�*�Q�Be���3ӏ
�e�ӱ*��7�m?6���?#���m|��>�3W �����նL��gmI�f?��kD�9Ց_�Bз�
�p;�r�L����Jmޭ�ܽ���D:���^����ʦje���M
������E���_w��})��� /���ou�.�Nx�#E{�^J2��šBb7� ���%`Oݒ�aM�8noZ�[3;�*����������h�����(L�Z�I��8�%l�����0��5�UNi�)���a���dm8�׏���`B-�YȨ�F/�%~�i~8xo"������Ƽ.�S�,d�A�_[��(\��EJa(��, ���?S�h���	��Q[�e���r9���-la5�>Zv�l�h|~#�����2�Y�f#��`f�`�:5���W����7z������5�`)'��M�A��s���l;*=�z37��z�a���(G��wR��W��f@��,�L� ���� vi��z����.�S��;:�J0Ð�ċqvJ[Ϻ��;�Mr��=��qچi�A��H}^y�Tk�*�K���޶��Ы�,�(��b�e��u�!*i�5q�����{b"��o�O�n~�w���X�*�c鏹2<G��۔�f�kf����w��|>r��i�	��Qe)�_�M��)�����*z#���h?C��Q��x�Q��#���J��+� ,y�`"�y\��ϱ��a8��k�~w�+s���	6}�k�<õ�f��F	~�8K��]��2ʼ�T)��]�|��s�O9�V�\�'�Q���Y@߈�!`��a�����!�!��m$C��'��V���ߕ���Ty�1M��pY�g��;z������E�~S&�])�DF����{�-�	f�C�>�3�
wk� ���o�F�v+��KX^�w��K�k�A�+������HЊ�˭Zm{���˙`�ZJ�ű�2Foe�r,�������])m6��2�?Iܳ>�9�G��"�%W~���t_�n�t7�IݛT���u砫G�4KL�/���Q��Z�!�×�v��TlX����H�ŗ/��H�$�D!�f�����Cr7��a��>��75ϓ09����;��"��9�C��%���0MT"�DA�� �ED�1�z UE��MǤ����쥯S�90��vbK;�Ǻ�to_F�!����bݛ�0D�I{��
u@�:��E��J�>)��|a�N�j�-��;w�U��\����Kv[f�ڗ�9c�*Jd}�C�����($ɌGp3*���7c�\���G�8t�{�=n�~A�pAێ�r�b!�|a�M���(����=�:$ds �h���Vl�*��ʖ/s���4��{6��$AQEH�jh�@ci}��b�6���3�d$�>$�*t�����<�~
��<<���:F63����B]����̳6�~F��cj���ӌ�9�ت�y�[��P/P-�3����:���o�*�sؠ����j��ɭ�;2�N���F�jVPwG@!v��f�x A�2R�ӗ��GDj�~��pg�d�6v8���?Ѳl�s�{Y����r�ڡ�1/:�q�1��H�敎;G5��Y�����װ+���� .G3Q4Z�m��X���l��W��r@����-3r\Ÿ�Gi��eXD�����N�<�@pIe{�|�C��1$���o{{Kn2c҈�������@�t�)�hw���}_N�3��Y.KkOo�c/�!$�,����G9�y�x�u�����8\��aZ���1�r�e)A�N����{y�lf��Y�d�Q]��:0�p�9N�4�3J%~`���f���h I�5�C� �_��Y}?����u����}{���ͧ�:��-�
kZ��}㛢Du1m:cp�G&��FU��O9���E�41�g<�0%��-�"\�O}��TO��T�m,�ID����)������\Y<�p���)��xԶ��9vy)R�n����C�z)XZ��{�R���(��
��ȹK��X�a��j����	��(��U�����Sݣ$�_M>5DV �&E�a�oj��=K,%���A����,����ـƷJ�l8�hj$��ϴQ�|���`X�Ğ���Y;�����0b	=lnHDȱ���R�4���Ki� \V�b�5֏�ذ��(��֜	�c�c��e��k]�l�%P�Z�;�0���OCO�x�]��w�k6����Ž@u=|��aE�Ov�ԥHx~׈�P$�
���i'A7�O���,s�E�O�
h����&�(x�hS�2��ҟ<7�-�܃��,��M6%jC�$@q��A�����󺇼[,���Ѡ�Ͼo��T&��#k�vX��l��>	a�RQHJP�Ӗx��S迆�i�k��t��.��(;�n���W��XU�%\�a�F
�^�"�͇���%Br�M�]�c:S%��,9�Y7�r��<��~2t(�� Q��:�����L����T���µ�"$���ӌF�I�sT@U��a3ȭ"�+o���9��z&�l�C�]�ފ�O�C�a�.=��_�3���.�3;@5�<*:v��h��$� ��Jh�H����r�;��:�:���<L?�Fd��V�+�H!m��<�Bx�9Ug��(�}�3G���,���#�n�����p�*���b����5�S�������?���;�q��V�A�Tq�������!%�����y��	�Nm�Q�V
��7���GHD� �!����Y�~�p�eV��H;lUhOe����߰.~�Q�
��4�(B/���=�����}����ad�|�C�B,�E�&u
����a�}�rB7ĬO{qNKu�W�D���?E
��o�e' Kڻ���d���k׫W�;R\���j2��%Tw1�7��?@d��s	�������o&v��@�<1]�v�31;l��ui�Rn'A�!��\iG�L���L��&I����N\�S��c�]Nr��(�Z&~�\v�=����U	��r��JS���qF���qw�B�+��j�1�^@LtEr�tמo�Չ�#�a̫�j��ο'���gQ��DP�L����Z%C�U>�qf3^�Nf=���&�v;������W3�8��k��2�#�s���tM�z&�����8���Wg������! 8Cs=����w��)�ل���Mշ��Ժ���@��TO��q�v9��o>���M������z�&$�p'�.W�*hEژ�?������󋾥�4˃&UZ�'�,���y!�����ɛ���qp4]"�����=R��\nƎ,`j�¾؍�Fۥӟ�gR P��Evn��E�x�$s�ۮ��sP����d?B�䈒ێ`m�-u��bܵ��>��P"�j���z�P���5B��#_�ݵ\Z�z�̇!���`ُ��y�WB��z�?5�T�t� Jj�Z����ȏ�����6��$<� '�miF`�*��ʜ��NAk�&./g�{!*�wDW���i=~��8;�u �L
�Cz�D���K�B��5���'즾P��i�]�CPw��[���0�T����^�$�P�6�u�f��1j�AԄE��E̋oU]zz3��&��8%� ����x7O�?L\81޼�~j[�%0Z%}�s�:q����I�Ͽ��/�3������jة?ޖ�-hu	��^s[0��&D�v�p�{��i�"	x��h�|�`�^��aC~{�p���VY�c�RY�T���cb0�0��[nS�A7�����'�ָ9l��sP�JK�v����3��~��ԈJ���W��V1�P_��C�e �;��w�h�$�����l��ٯ_$"�d�Ê�{`��WDK9������l�N��aEg����>�T'���9Xht~b����59�"��G�F�BG��L ����0�f �����#�9��be�yh$J����\u.�R) I'Epm\��A��P.z.��[������Dп�������TdH2�z���x{���+h�Ԩ����]�}TB�9A�ώ�X=ۡ^b/B�ڈ�y8f�N�Ev�b.z���������b�s�����y{K΍|��O.f�y/I�@m��_{j�"-�)V.�{4pB �ӈ�si�§UOƘ���#��]|�?�y��!�c�@��Ur�l�~�'}1&j��/�ȋ�C��G�	��Ehd�jEg<�&]��/G�O40=�����H!�	�p����j<x��\�9�T�:�T��%�����	3i�N����ܥ�Z�5�����cq'��A{/\�z]��5��).8�JPF��;huD�5~�<���Q�D�g��^k���P�7/�ڈJ�Rz+ ͽOy��J ���/f�.��;�����JͼX�y�h\IE��>d��@�Ŏ��������$��C�(鐂qIԪ2Z���|�I�p�6v���8��@s�_C8�qȷ��oCl��Z�jK��L������D����/`�X�$����K�B�Г�$�i��\/5%�5�f�G�X�}9����I�V��XOX�Q�j%����Di �=���b����F���ڲ�jV��@Sec����-����)4pmoQi
��+��f�J�$[��6���m�S7}a��f̺^�;q>��8�f2�k^E*G g�g/�@y�fpfK��!x���*�����a�+�f�8"���.�����{�SH{�����cRZ��
"������ZьR�Y_���^I]g.�����v�ŀ:ّ,�&���mt� ��7n�gC� l���|��y��A�#_c�tXFDjn�	b9�w��Ǐ /��:ACÆ��ے�����Q=�WD=�SF��m2�BNF��(�q��
P��|� �m��,����J�6F _(&�jM�ᲺF����O�Ec"(���r��q���s��b��
�P����On>�B���c]3Էܕ�L�3H����$�iܵ! �7`jd���bj	s��OK��Ninz�QM.��63�|5�(\��@>�{�,�o������ݾ�6����EH<�g�=���1|z��A������	��'�]zC���n��{[��S�"=��G'��r6�˲a�]%I"�Pc/���.��{7�VŸ�x�Z�O��n������D�me��07� {<��׉���A_���#*�D��c����[T��<���b���  ~�KVC���	�;b�!+�s}e�ӈ�j����5�M���i����陠��8�pm��=wü���ş{K��\��X��֑n���R�`3�f��2�~���M���Ɩ�{�b8 ��BR�'η��dv����j����|��/]b�&`��V�80�ʿy<D�:�(�����QgĿ>�w~�A�Z�g}�=yCN&��s�K���X��S��JT:B�� �aq���7��`�6�5d�S�a ػ����jdM�7-51
n��X`�Ú������#QD��	Y��#כ-�2B���2�c���QT�g���l��x-������8k�#�d��5�JD	�-�Y*%v�۞�በ�����Z����n�P����n�ϥ�1�x5�&�AM����2uΤ�V����nAd������N��4�5�����xߵɝ���
a��i�h�0�P�-voE���
�o�&��Oēmt��^9Ҁ��7������Y�CH,�v�M����_�$�kq�Z��)��/���(,�q�!2����؝b�1y�w������>P��˳s�J��f�7�������^k��1��L1�޹����������K�X(v%=Q�GM����W	��n��Nv�rjf|�:426���z �r�l#�-W~����^��;�:lM����L&��U]�N.F�U��lʌ\�T�VB�aT�v"�zU�@J09V�1&y 6�k�O�?�aê˦2`93�+���;��H<�rl�kG&��� �����H�{���;����ԣ��D�L@�G� V
��Hn��m:���>39�����~@�h���m�e\��^�ap��f��Aq�ב����S؉g��.���ܚ��}S�A��q��$�8��-��������ݎ��]mb�V둸�8,��h*d��ᛂ��<Щ�����1V�p;m$�hp�·���=�QhL���Pr(�������R�}���,�#�ݦ�Ֆ�YB��[���P
��C��V�}ŧBx�O��rN�CW��y؞1�
��#o�˗AqW��m�d]M���U�W��G\d:1�K��&+j1?����Dd�	tz�K��0z辆��A�1~!vG�;�~�8ֵ��F�'�%E�]"��m�������i�L��ߐ��]/t��������&�����\=c��&4	b�1r�_9S��m�AP���P��1���ɿҔ�@�Nr΄Kן{���
#-������󴿿�~ĺ�Ro�nP�����ZR�L̶'q�{�^]�=ot@&�(%���ҙQ�y#jk�t꤯�s}ʍtwO&��i�+�8���W��V��4!�/sޚ(��S4�
����ŘM5�������8E�����=qX�eڡ컿wM�4��+�����]'�8��륎�yڎ?��b��y���4,��U�$*'Y.�,�V�yM����H�7�Y#4��ه����}ǥ-����VL��F>O� (�R�����ܤl��Yxes����o�2��Ű��e&}�/jM`.�-V�����=�3K���(�L�yz)�sپh_Bզ"#`��}!�z7�������9�(��:�B�}T�@��T�[4�A�5������ۏb"x���t�i� (^�igI�*7�ʜ5�PA�4_.��<� ����W��zi^��.Ѝ;`���\CC��D�1�,�~���N!�'-�P��LC�*�払ЌT���0�^EP�^�uh����.A��Q�x�c�p����j����}�=Ɩ�6�Ex��� �9/��<�[��&���%����W��]��Iyⶈ	�T�������&�1%�uʟ�^T�x����3V��y��/�]"�p��	�2�!�^pA�C�<pÂ���������Y>>��"}�0{~K�<t��B�%�����h6~��zp��*xJ�C�ہ/����𱺅(g<J<��W!��V���_8���&��,�w��$,ǆ���l*�[�Zl�_�n�dt�|�\Y��XY89����]Wlt�n�8�����h��Y'�7�9y��~��aoUc���C����;�#�䫟Cq���_�qp� ���R��� �IvJe�e_$K������.+�� ��E��6�u�����z��[����% K��a���վ�<ǩ�aH��z�w��yŜ���+����	-U�&+����G�m|X��!UbV��;�by�T�fD�E7/b.[<~��$N�.0>���sU�R2n{�
|^]g.G�~0�F@���_�����6�)�c�{�U� �mY��DM�õkUp���]ӈ)�n�]�Co6zy��6���A3�U���'�(�&�/����>3�b��G����fXv��9�<Y�t]c�/��.4�:��s���I��	����@�<s�#��Д����F�/���l	T{�N�B��=�)Z_ ��R��$ ��{�{0Tب� ��v�>����+>�V/h65_�1���ݽej����nb:����{��N�Jf[�+%I�p>���i��W����������R�J�[�zI�\,�E�Yo��0�cM�!<%�W���.(ꗂqj��2��+���Ir�6E>d�|�!o�_D�@q�/����C����AK��jL[r���4��- �/���X���/��KH�Z�Tڱ�JK�\��%�Ϲf&�Xx_�}��0�BIUm
�9>.�Rb�%�#������/����S����@�Բi���T��axc ��H��-,����.��QJ�����2هd�eL�2P%�v�Ǟ�H�}"2�f����<�����X�o��H*�6U�6ҴT!fQKwK�Yx�A�;~���k�aF���}X8�`��8���č�{6ΔL�GV�B|fR�*���^�}^����{b�R�_V�^�Rg����`���(;�>,I��R>�t�.��hGg��_lt0W�]e�z��A�x�z�t�E��Y4����PG�ΨW�/��EAdU&��^�<cے$���GEE�4_�Ѣ=�c#��Ed2(AU�H��{X&����mq��,Jo��.6�*(���Mo�������??�0\�c#?������L��}`Ɯp��p��PmU�0zo�CW�� 3D��������X�mv��*��!��`k]v�1jJ�&ܰ0(�ϣ&nD�M�_6@)�}�Y�I��,�{�����K�鄞�%6��~�H1w�g�1��1����$�P�լi���sL]����_ې6�r���"��B���S׀˳�]FlS"R�/��.!�V7�\��I�;��O����4�G�=Dv��e!<F7g79<Q�X���.���~� 1�d�]D�:�#1���{u��Ϛ������2���V���jh�b-J������u�K�[��E԰n$#Ϫ���?���!'�m��p.-�=X�!������7����U��cĊw���OjR�o�3����Sw%�Ͼ̗�*�w���� ZݕR��|��Sd��ꕹ�ey�����م��p9�7�-0�Zy])r:ﱿ��f�Q�>N�|�7;�g~��yd�(���9K*�5���]SN��T������b���47D`牚�#�S���|��sָdNyI-V�Nn�P0`��e��A�IQ���� �$�A-�[��x�8l2	�������"���m��$X� U��F���a1R�"@�%�]9�
&��0U��\�O��a��3���3 $N�lx�;>�m<�+�%��)#� ��p&[�H%�]�#;�t���n��eo*L}0�bf�V���H���m�E��@+�9�g��D�a����E���?��c5�D�W�[#p���d��/_��USU���:�>}��9��z%�A5�{�C6q��$n��;��ʡ�k�	hm_��V��u^;�E���������*�W\�.F�V�;�C�hM��`���o�Q%��}i( ���`����^X}�a:���������S��B*3e��l�
(.��P3}���B�9�O���N�RQW��Q؛d�
0o+o4����G��dz昅��W�ޫ\a ����c��1��qmd<G	̝"��}<�-B�#Y~ԃ1[�)vģ]�B؂�lV�1���H�������9�J�9�
����_�	 fZ�U�� ]�:��hD弦�&<ۤڹk= R۪��	_!�r{s�S�?j�o�ݪo����ն=|�/*@
��rk�������#� k�)\��E>Y�~�ķ�4��P��י�V�Zϊ?��[\qP3�^�ì=l�&/#���_������k.���a�Usچ�t��&���f>8�l�W%�t��!^��s;d���H�ŧ�����M�`�>ԃ�)�)�\�\Mg�qU%��>����M��Z���5Vbɒ'�¨���	�?�������|ax4I�ZUR��'�%,~R�y�ȱ���`��L�4���D̷�;{w��܎��I��2���F�u���R>�3�C�ܡ�����s˩��	��� ��L��"F
ی�~`+G-�;�쾎L�׌����N��J	,�z�� ٻ�BrV�#��ݵZ,�z�ׇ������?�7|�B2zL�}�T���9R�ؗo���j��`����xᢲY e�iDn�*����R�kA��.-D9�����W7[}i;9T����;}�����Cu�D�u{�ɡ�8��_�'�01P*l-�VN�CN�x����� �T��n�^���P�u%���/�LA��V�4 ��x �~l��")��M���3x�r����vM���"�[qI؝Z%����8��Z��I�L�Eb�1`z�N��:�ҩ}�����u�d$^�#����s�V.u�LA"G?u�fN�xe^�?C��6p�ӏت�� �Y�yd�00x����rw��ۅ�&���Nݱ�JIp���M)/[�-qɅ#J�+}W>��Vo�w_��F�#)"�Ēw޸�$	� Ó0�lGiR��_"I�dq���>���9�k��X::l�����D�_���Ū/Ƽ)�'8�h9V��~ �#��f�s4� �Jj���!�ܶ�͸���O 	��ix!��F��eu2�$�U���,�.�"� ���E�$�����ϑz��[:�����c�0�5e�S�7�
HTz$�߶�E���+&���&�M��;	�{/\��{�M!�XVj�\0�bӘ�X*�yvҮf�GOE4�.�<F��8��悪s;!6�p{I�I|[�.�͗m�@k��_9=���
�)���{2�, ���̀ߴ� ��UMJq���F�,�I�̒$y��,����~UpU�~`�'���&�>�/�9��������G����C(�(�<v�] <e/E784�|7�A���7	�NHʽ~Z<����܇�R�I�5�����	1eNUh��Z�|Z������!��w��{m�ݨxw`��:��b���㳹Ph3M`5�0��-��B��|�O�5�m��!�5&$�K�J�+O�w�Mϔ�'�t�ώl�E�9��O�JJKɯ���\	�>��2��5���̏�~ �Tm|�C>�('�MqGf�2�Ԥ7��I/��6t�a����_��Eq�g-����C��HyK�xLX��z���J���+/@XjY��
�K�ߛ�Q1���\A��%�!f��wX���}C���;=IRqZ���~��Y_%�v��.��9���E�����=|s�{�8��>{cc}�He�5-����'++��Q��7���d���`O���3��h�}=�fJt�yM���s�JJ��*�˕�eb%���f�GK��x�ݗ�����a�G��L8���C� �	t��}2��}�daf���*RXqN��p����?��X�bRm׬_s�^E.Ag,=��2�8x-B,�N��3�t���u�gAW�lq�H��P"��D�A��)tַ���+`�M`��E�/���AA)�l�?Y������O$t���M���@�$���*(^]�h	��a��7�mZ#,Bp�h6Ԅ(��JM,���i��_9��{;c`R���I�G#dǚ���Y����K,Pj"�����c���3�G��`��q����$x�'u!~��`�J)���(j��I��p�����nx��M��p6�F_��yP�&(�����{8����3��g�����6%d;�E�H&og=�ɐ%j�1�̓��M���I
˔�'�]xK��fo�S{}��B%";�ށ��ē��]#5�"�6�/2/�.��7�KS��$���0�O��3�~�n�Ē�D��eޠU7�35<N	ԉqY�\�]^���&D5�+����Y������ʟ�y�|�V}v�Cb�
�q�1쑷s�� ���ҰK!��'��\*���ҍ�ʥsp+��=�g��;ŝ��9R��r��{���E�ˋ^R�+3����0�~�L�H�9%���:�`�p WƐRTշ�ondt�g�ʬ���ͺ��-$;�����	_0��y:ZO:l�B�C�Q��>�\5y�Vػg���yA���s'KG<Wʖ��S��T������{4��7��B` ns]6S�-�y=֥dd�I\-3��n{$8`+h�Q�e���Q	���O��a��-��j�v3������6�VR@�u�s�?:���kyO\�d�5^Q��볳Y�W�!q�jk�f�T�/�ك�l%R�g�n��w��iw�v�&V)��vz�2��<�Tz���!~n��mS�� ����L�a��wiwKq�}1�@8�����̃�8�B�-.��kM�=(�ZWV���^"��BM���l�Z]�g�%�f��o�tI�h�"�߸�0�4�V9�� �|�F��yoP)\ta������ �IE��
ѹ|k�!~)l����G־f�7|�1I����"����?5m#n�$�2����0_��k����0�k3��<�#Q��f�~u�� 4�ذ���>P�0qp�U��A�@uC!��'��O�k�����1���m����O�ׄ�AX���f��:i&����;�if���	��K�	~��G�|)�K�h��r7�r��m�2OI���kv?�U�G�>Z`ڟ��.�1P3�j���%G< ы�-ǌ�I�>V��#!��P��o1u���A�9�����N>�%Ŝę�e�����gИP��f�*�w�E���1l��RO�eư�*�&s7��6��?�q��p"�l�W�]T�@��P*�L��?m�K;?34�D�ϑ�1x�z>�4R���L����_��Ph��FY�eGX��i�'�^�{���j��������4x�IJ�����'0�Kݪ �ܡ$�z��e�x}`E�E6�t����ץ �K�%��cח�;�Z���;��2��������J�(o �wz(O&�ZMgL����lϓ�#����L�՘A�����d���U58{���jkB�
���-Y/�F�6�%�����o唜���Z�?�S��q҄�[Z�\�/�����Q� �Z�?֌�h�M�	�e�[#���;-�)Ԛl�-k5��vW��h_a܍O�`��ZDY��E�(�ˣ#�S5�Z������
���������
�h��'����dP�se1�O��=k��D��<aY�z��O�y��	0I�\�o���G��ßv�]n�=tB�s�.R2C��o:����3��Ď�Iv���[�/��9H���#�� �q����H��o���@}����9~tЎ�/�k�bF?��x��*̱�4H����ab�ܒo���n�a�w*�?�["@*��o�|�d<j����N��h�wO��|A&���̂AQ�Hu�P�06�)DY�%���-���'�?ϕQ�&{��`�#á����t+}��,���ê��B`Q���C;B+8دi���+w԰޶[}��<��%�ƱF���8.�|]���_%{)��U�߃�s�\�\jP��V�4���5'�+=�`�?ϒ����0�߅�C:=��^�~�8[��W)1�0p�夨z���夑��9~��>],��F��>E��,d���F��F�
��7�6X	��<Fw��+c�X$�ww�����A�-���_^��"�O?���m�qX�No�=�z���2��u��bhۤ�rmY��2�P/?,��>bFG����(�
�Z��_� ��>����T���u*\�G�X}L�� ������r!� ���s�TOj+�<��7_yŚ�.�T�v�!��	f)�;�/rrV�-�_k��A49��3���������_�{�gĩZ�Y�����7M�����#&>�G���-a㍚�u���bV Ch����L��5᧓Φn��~�07�b6V��z.t���ص��G�f�2�[w��Կ���u@Χ��wJ��v��d|aaRN���-y6��+}w�+�������[��+�b�!c�-d��.����_(ϻG
*p�sAODxcJE��K-�2�t�_�=�q~#d�p�_"�=�fL a2��ʹ�R�՞�=���/b�k΀3pМ�����ʁ��/����?{A}�$�K<E��W�;�`i��;��((�d�>Ux$.t���Vu�
\�Ǳ'~��߇�~�{6>���`S}Bߓ��6&�>S�~12�cd�)�L�*�D���u|y�t�;��P�&V$��G|{�~+��5���v���� j%L��8��2�r�!���ij)v�w�a�vgl��� �n@2=�y��^�Db��#y}����/�c>��Nѝ���NY���	�X�E9�1�����U��,����G���Y�7����e+`�ܪ�M�3|-L4�9���L�D���9	ߩ�@����3�p��F�ąy0'D�T��N��;@ۑ�eF*F�n��1��z��7�{Ǝ3���ғ��ijM��p��3Xh	g�h�s�~
଺��Kvl�z!�����Wܞ�W�r9�u�x> 6�H.̂CTZ��SЙn*ӆ���e�FHN|C'����Ed���({�e���/�N���3���`��f���T�FI�?*�n�� EL�D���H��u�֯����S?�r":(�*������{���u��:nԓG���F o�Ody���"g��u��8��\��}��fO��pT:��4�n�.��)F�����\�c�S9R��_�R�ƶ��p�J�)�(n��#���`z����`Z�ծ�����U�L�dƱ�cg`zC�����I��t~U�1�5��N��7�Y[5�Qc��;j���Kw���y����^(�(\������u�8�"j�����d|U��k�r�	��$�����4�	(,6H��q��]xRq��+	Fi���V�&�5a��+#	��R��֧ hc�[2�0��k��?lx�C�����0�XONA�xS����ka��𑍮�+fF|	 �Et'��rlx�E&�`�
뉙i��@�:8*�w�yE���
sP�0�U��{�Ҡ��Ҋ��7�qh�J�<�SM,���M��D��$��q��n�_����K�,�p�k���A�ߑ���d������>B�˽�lJ��w��M�ޮ���:k&�r�O䋷�B~����9ڼӂ��X��%G���ȭ	���!���x�V�&r������:>3N���l�r�I���<~��F����lY:v��@��L�Y�d۔X�M6�w�ѷa�^�^���a��|"��#�J��9�zO&��i���O�_�aMԵ���h3�@F��2�;k��<�" �u�/�6\& m	�s/H���=��;^N��}��W(L�&��V�<0HxNcm�z��m�:9�����Ã�^=��7��W����I��pj$��(9	�V����S���'GG
�8�f!u�G�A�:�Pc*ɛ�L��������DW��4f8m,�V�L�H#��ϷO+������㣄X���LV��;��(h�g��;����Q�'p���(͔���T����}�GS���İ窂��d�BW'����}
���q5}OBB��O�@�N2gW�#�h[�
�?�oA�v˾��l\dg%��6/�W ��\.�h�Uz@�p��1��N��5d)� 	Y��������I�,u15Fv3��q�����8���㣧�T�����Ws!�&��������k�]9p�:��i��&�d�l�=�b���	,��r��|S���!E���ᷭ�۶��ѿ\)�@ױr�c��;��߂#��T�I���Ȱ�IZ�Ą �y7P�ۙf�1Zj����q���^�|�=9�&��J��������Cr�k����؂s�t�@& �n�D8eQ�WrR(���!�*shו�y!I�w3�.M��K�4���z�;q"{(ګ�	�MZ������3U�q'Ix��ǉڃ5�?C������
46R;U���'�(�,K��y�(�tNc��y�4�+�����hb4��6�'���f���F�R�
�iR�!�p��n��c9sؚS�B���x��ϾK����۹"v`��2-`�S��<E�������*�ՠ�� z�Q�و\�B��#������zw���}K��1�/�'=#B�T���EyT;h������[VO��e����� r��i��*�y�?g�A6�H.ZY$Y%���WD��i����;jӺ~�CJgDu�g�6ӈ������'���P����k?C{_X��\�O�T�8�^���PS@u�C�\MkA_�J���z����%���˼��|�������x±��*a���s�@z�[���ŔD%H���eJ��'�}I���Rd���/��'8��
�f�� u�v^^���ѽg`{�e�9r�"ԍǫ�n��띅^z�dC�~�pM~��aӸ��Y����-�0E@�Fo��,k�_��2͋���0�>�FJvJ੥m_�H#�:����6WJj6W+��V��y_�P���Ż&�_w�W$����k;l4��1i_Oݺd>��f���Y9<Nf��r8l~>rOk�����ݒA��)�9'E<u9<H~mHym� �M7)�}X�-������zU�;�F �&���bN-ݘ4{e�ܧ$�M�t&.�QF �<E;[����&\�yz��[+�	�Ks��տ"?��S��3�xH��z�����q����S+s�C���p�Ǩ��ă��"MXcNg�	A'b ��E;y��f��4E�G.e[��$$��9����Ss(���G{va>|(�.Q	�z�@ƍ_�]���4)!#�{_�� R'U��7��
=U�q��'K�3Jح������y���szË1�U�"�zv'��&5 /M���Lm�lWBG����	 �uw<c�0]�ZS/r'�4�r'�}������	G���
��<}k8�'8>�c˭ߧ���8�iZ	� �N�y+�G�`Z�1��������{z�L�%p��@Iv������@h �95i 7�����f��ɡ|�"R<��b�c��JJp4vP@}s�K¾�l>��(]��8F�&������6/���
��Փ�e��XF��+��X<�w`����iA����"J�x�}�ր�p�m��k��'�����+�2T��@���?��/�mD�2Րq?��i>%�G,,��	����&_H��ܞ�G�THP�u5��G��#L�К�.��gf�!�Y��D�hT����GF��5��e�ʮY��r9!��)ft^�\��ra
:��|Q�s���K�~!E��w�ߪAB�r�e���3f΀���M��������&�h_�-l��M���f{gb�-C�;�ձ$��'�><Цy�M����0�ba_ǐ�%t��2���c�q��t���j���@�W~��pJ/��1��al��NT��-D|X+>w����p��F�:[|�^�mߧcd�ydӼ�Y��~�u(���GeX�pI�oZQic���dǕ�]�tz�%=p�~n�1pW�H�m�	�a�>���֫`��=��8z�C܆>3�;����EUʬl)/I_O��n{��$W�E� �d��i%�8�8���Ҳ�+$�w�� п�u�����~ �]��$�l�6�Z(���B���m��	�f~\mc�6�7;���v���n�y���˦�LP�D�I����8��iy��ض�;����j����^�2�D��8ǥ���jt�
w]Q$vrQ$��� o�!2h���q�.D &��n�)��.7�:\%�Z�������GI|�Y�+}T�*���1Zr���P�q櫦~G�[Y�q�; I+./��Ê3�d�4�^��ϫ��ς��$�*<�@��]�9#3㵸�j���D��?llNQ@��weQVm��F�1z����{Q���I����}�<���\�-�h��p��O��	�>����K�Oc�%n�Ǐ���v�"UO9� x��y�3���RX�w��y�I��LerbN�膯sZl� #^}�zO53U�П͜���N�F�3 zu`���4I����<Iײכل� }"�oE8��Ƕu��e��U+�ŋ��}a�:���`~J�pp�q�u�Ȏ:�>`G<<.F+�kO�ôЛ�U/e4gh������|�\53}��hOLF�T�l�_.h���)1�3�8��\o�^q�yJZ�n�XL��)�n�qn�Y�z�u�*\M>,�ߛ���O��=��鱋�ֈ~x�U���|X��9��X�mutO5`6������Oj�rK*/�d�?�k4��񇮯 ���<R8�5�j:hϊ̙|@����?Ĵ�/1^�E�O���A	S�FH����]RS��֔�i���V[I�5,I���Ñ=�`��}xc�bN�;��k�9xlCՇ����d0�s�O��Lx����k�<��\3
�V�|�DeE_��*lx�B�&�
V]�i}��e�г<�Er3~
��<����lxb'\��p�ҵ�B7sl��5!��X�,���M��7�$��
q�"��N��{R�����,�QV�v���������9?O�L�?�d[>eA��h��J����,ًԩ[��G&k���:a���\d�!ƁD����X�M�%r)O�,������l��#����r_Қѳ�j:io�s����^xr�|R��~|�S#Q��}:��f���5L���j�O���X�$��"䌜�`ى
A+0�a�[�"�1H���y9���&n�L�^����Ou2�a8��G\(3���S�;�ٱ<�q������� X����tH����H�h;���ig#��zVL�����V�H#�m�P��؈?9Zx��ܩK�SB��ڂܵ�9�7��Ο��op5Dr��A��ަ�p�HS������K��.��f�A�N����iɆ��B���먡O�����\m�VhV \I�=}��UP�nS�7h��C����ƶ,V��;B:�h娕�����D��Q�D�Sf(� )��Y�}m�}oCX�Ai��M���\xB� J�p
��[�v�}:�B�fkO�^�N!�W�϶�3�
�:�o����0����d���A��W��(\��@��p$��T(1�	��4d��	d�3�@�i������C�1��v\�GJ킍gyo}�g�7���2V��BL�sJ<o��2Y����6]df,V/�T�&��r�=�|��:�	�Qvr�Sd���:��߷X���վ6�ǿ�@��rAS�t���k��#B�����2�ݘ���+2�O�o�6P��m�Q�Zgw��k�Cq襷^R�r=�9&Ǯ@���^�x�fގ�<k�Q���^bsrd�t�O&+�n�}>8PV�W��Ԁ��I!�c�s�Y��D���?@���M����#������O��t�q����ɂ��a�ME��������'yAx��͈ڮ��?������]4��U��'N\,Cwy7�%��'U_?��!��4s��ε���5���e�B���v�wng�F1� ӵ�R�����*��9�s���scP��-�ܿG���z���x*�$�`�H>-����VM��oT�HI����v�zq��Si#B
�f#5XF���<zL�χ7A���<�������B�����T&��V.J�pf�fj2�W.��LV	�:F� ��i�G�*L��� �AA�X.�)2�6��-7jW�y�i�*�C�;Q��"H�C�r�D@&j�ae�ۣn{i�'Bm�P�;Z���C�ȱ��F�bT94���^+��P�}su������A*|��'I�Ezv:q�ِ�N"r�@,�+y�x���U�L��+t�[	΅p�%S����A���ؘI�z�ݧ3���~��_`�ӗ����&4�u_��^�_
���^Ѩ�_�)S��~"�yū��J����^�F�CTx�p8�珬�R�y`}Y��1�֖0�i�q�n����Jʦ�}p��O���I>�J�-�p�B��p��g���קJQ(�W�X�VH_-o�໱�Q`^wv�"$��A�+E�l�2���|_�69d	kX���+�- 9'e���f.l)�&Z�������]c�T��'��a9��~�(g$f����K�:��Xg�t@�e���z �����K��7a�ދ�e.X$ ���_n".@�x _��EF��j.'ГzD��[��k�N��~�̈́���MǞv�HZ�9z�	��N�ӌ��+�35Ծѱ�{f����̏�:�dVX�՘����bkU���yyf9ݯE�X!.��"�x~��mj��sӈ��w�{�R|�K�.|A���@��_�)��8�j),.�{�ju !�kE���hU�S�r����ɭ���dpEyMQi�7�i�%�U?�}V'5F�&@��/�/�h|�◀fG��.��)ӓ�9�<�K]���/�D�4�=� �~x	2h^�U�3<(���2���껂��P�;�'��m-	ɖN������Z��y�z �乌���I{Zu���ǋ�4�?ϡ� ��K�h�U�5�5�9��rG�+>��/���͓�����J�D�+�4���H날�L�=������9u��$J�d�O^/\�N��2����v�d�>��E����ۡ�(��Yq�f2�h0���hI��6�G�!��V�q_Ϫq^)0�/�-C���0�cK�O�L�����uQ2��B/�LX�	����6K=�5����-�\ٱ�%@�f'ؘX-T�}�6��8�I�!,�n���'�_%3}���S	��8���5���Dز�Vx���֜Fc���g-��f��Xh��kQ�������PO�z�A����}����}�5)f�&����c�5��櫁ц*�ֳ������f�&�KVT�x{�P�����BaYj���,�8x}���ġ";��uΩ�1�����%�R��(�`���k���Ӎ�(zR��_Kr^݀1g��7�3x8��r�,|���g~t�K�	g�Xl	S���z�O;KA�ˈ���tnG)@�J� c���8��+,/z�A�
&����I��y\��_��I�i�������}|�Z�(�ޙɝ�p�̠v�am�%f,ڮ��Z��6�+(<��M�g溩�yG0 �e_�c����?Ѻ���2����Q�e�_PX�e�����53*��ܫg;�	���br�ԿZ!�c`@�P��Aj_mm�e�F�$�ne�M��86Ir*�R������.�{�'��E�A�@�V�3�;6���g�qH��wg�x㐽�(1RNH���}��'��eꔂ��]�!���g��␵`��"�o��>��8�ˈ��]��0"*#G/ʮ�.v\�7w�@�	�p�hO��x��S�\�AD+�Jev+�7\�<��	�,ȠrB��f�y�LD�n�x����z����;�$�������V����b�C��	�M�)x���k�����:Ͽk"��	F�v��b�/pÔ!=�S�����5�Ѷ��
mf��lZ9�c|�R/ 3�o�����-���'�j�~��5 ���R�#�y��d���I��{�R��őg�|'R�l=]0q�zy�Ө:�ˬ��lQ=4�>C�a�pjgSR�y�I��cKߓ��.�SC��T��<��7R���7�`�o�S�8"��a���\d#8d-�b�n�`����bs�u�Q��غ㿛���-F���@�Hh���E!�% �@-�׸ �0�qq�kt�z�5�q����dhY@;��W�tu��T,�k�qF(�;���oTn+���{���?v&�}6�b�2Kxλ�s�f�nW�<SH�̀��Q��gȳ�Fi> �wS@ж�4���rD��ۨ�Ų�ș����2WZ��@�"����㭕3֕Z��Hg0U.f��noK��"3���4G�ӓ��|I�ݝ[��o趹t�����6� b��I�m�
i�q|���!|6%5�]�O�V�7z\I�3�@��}�ן�#�$�> �j�S��U��;5.�j0;��у�~#'���f�u/mr4��5�E��>�#�0	AU2v\��b�!W�S�v�k*�$��+�³�'χw���<� 0X�`8���o�ҧe����;��o䈥;���ס����lF)7/�h�ꕱ
a)rC�]��>E�*u�v�@ZU,0>�[��7��ɑ��(��Np��{ŌcJ}>�R#�(�P9f�o�:�2aP9h�d���,�V�ݚPӜ\8�e+j�z�����M*2�͉����ɯ���De^:�*.��7Oo�6�-v?^�P[�9��W{,B����?L8m$��?���D6x��Z���%s��ڍ�sLbh����-e�j�����n��QO��^5���<�j@)(�w��z�����ո�<���3 �\���L��i[�x�%�Eva��̀��}n 8[%;׵���6��X�Z���;(�͛�֒S����Ӟ�Aŧ�C(���Z�R뿓Nlg���F�WDc�0,ԧd)����"��8?8+�����BH���i��Y�1HFj�%�y�oo}#s�D
�ׯ\S,Ѹ��H[�T8\ PKE����� ��
?n9�hq�	��2[���)tͭ�Bl]��5F�Ov��Kh����4��4��Y:Ӏ��`q��ե5I��r�._hU�1j�5y� +�'����s�%��=��#n�3�Fa�䠃���2S5   *   �L#�靱I��!�d��8�L�:�.ħ�~��ק(R� e'�(���(H#b����o��m�uɘ�2�.QJ�t�p�ˤk���+�4Vԛ��t�8d��	�9��	���C ��.1御`th&k��"<qmn���B�I�%�j�؁��!U�5��S�[1H�>�RA4�!?���1��6MQf}�n�;$��@DcӒ&,,�P*C" :郬X��)��"�*���ƥ���H�_\ B!�8/�ԅ�@��@WXek�+م�O�$C��D��y�8u��!veό+Ӑ�ӓ�ҧ��T�n#<a��%�$�*��U��勗(/����g�55#�C��O�tP��?)���ԁA�"��������Dx�L\�'��5�'֘!��L�.b�ir@�z�p,�O:)Ӎ�dT���'ƈp;�m�?;?�8�D�-G�X#ݴ�N"<�5+��aY7f٥L�L�8�g'N��G�L��>"<�U�)?�3"˭�i!��ӡ"^�p�L�IyR��u�'J��?	V-���)"��6f�8�*E �N#<��C)�k���$߈u,����˙?N����'I�E
1OB�J��$V��ē>��d�K��zZ
�@# M�X�~P�'j�"<A�2��<�CJ:p�l	�e˲B�<��f�ޟ��V��z!lJ{~�3?���*��'N��7mHf�z��V!}k�{��T�'p~|�O>u���W2o:�	�S� 3���w[��Ёቍ�� XpI��L2և�MxT@铉7D�\�  �݀                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          �    T  �  �  '&  y'   �L#�靱I�8��tE*���"O�$��L�'bj�����΂<4��ش"O�Ȩ6���U8�	���*�)���o�� #��4h0�`Ü�b�ְP6�	;D֑#�����g� s��q��,I�A��Q*��;d�����g�z�g��D�tq��\�WOB��&)B�m�1���/L���4��{���93�N#7�e����~Y�A�(ۚ�賠�YX����*�$�N����,\��0��M&D�����, n�e���R���0Rqc0D��i��J2?�e���*���u�?D��e�Ӥ9HJ$���X��dbL"D���A�(s�ZvKP.�H`H!D�������z@��34̀S���p�#D��a�'[�8`�v�D�*�q�4D�����8O(�ҒOU�ra�0ѷj4D���5���F����%��!i���m1D��8t�M�rJ|����"c���)D��n��'ep`�W�S~(����6D�PZU�]Qg8-�j�#/N�d�5D��`�	֋q3�����n��4D��ڀ�S.��ԁi�)�ZD��7D�LⳄ�
�1��L��<�d��#D�hr��)_ �5!�''Ҡ)�g"D� 8�Ʌg�1���-G���xeN%D�<�`Q�91����+����b"D�@��;^s$�[Ѝ�24���d�<�գA�%c
`A��B
L���0��C�<`���J�S�)@��̩B��g�<���&'�n(dj��H�h�M_`�<���{�#�W�e���s�`�<!�g�BG��R�,�<Fjl�Y@�y�<!l�=k�R��#�=)�@��%�v�<���I'PѾ��F��/W�4q�E�s�<	A�	~�&xQ�	�Lr 9qQj�<�VJ�֭���$��XA"Cd�<���;Q@�1���E��d:�i�<�B��Pa��3�$2dt$�N�<�gg�
�L�!�	�0BԄ�A�@�<���U&�ԭ��mX
 #*���"\v�<a��7ۼ�蓫?U�(,�@ v�<���U�|�H��#j���SC�Pr�<v�*lj�+u�H0�Ri�X�<Y��94���1� �r8�"J�<���ʋq*t���4<�`�Y�"�E�<i�NB�Cy���5
�w�r .C�<)5�>q��S�c̙�m���D[�<�Q&�/ ��YD��<^P��siY�<�ӣ�`fH��FcU9EP�+�S�<a�Ԋ�Dѳ�E�z��)q'{�<����!eƮف��݂W%x����m�<��ʓ({�nPD ���T�`�<��M5�DȒ� z^��SE��<�4�ͽ^U�H ���<��]�5�Cz�<�w��i;i�ɟ>5�23�"	s�<Y���.D��3A��8����N�O�<d�أJ�(b���i���A��YM�<Q�H^Myޱ2�bZ	%B�32��O�<���%m�r�2���/b:Ղ���p�<�gύ�<�Nq2��O�L)��B�M�M�<u��V��M��`ˊ;_��0A@�b�<i�B�pb�MA(��4)H|��EX�<��MW��p2���y��U�<�#�+9��� $ڋ5N��F&{�<Q%�U�?@V#J�A�H�jD��u�<a�fR1]�L�QN�QJ-���y�<�lG�=	��r�lV�f��BOPx�<� ���Ec�b�pyy�m׍J�����"O�@�V@ό#+���"�WG���"O�T�`�ۊ�Jp�p-I_�����"O(�A��:��	q�R'K(��"O�M:˙�d���Bu����"O^��l� %N5	"�m��(��"O Y�B�E##��r ���R~ԁC�"O��G�Z�.�^�����8Met0�"O�Yy`E>J-��d'F(�"O4�B��B��ݻ��W�1���Zv"O�,���K,o��ٸ�I��h�,�3v"O�$I�krQ�"*�K6��"O�j��B�L�����;7"H�[�"O ��X~C�鉷��'f��!�"O��
�b��=(��\�C&"O(���c�\�5��I�'J��4"O��q&b,�Ŋ��^���R"Of%bY5�v��6%��e���`"O|���ف+����a��3�`4��"O(� ���)/�a� 3�����"O����ѹ0���⧞�n��d��"Ot=㱪�t���+� E�*vmش"O���g	�;{�0���G�*Wb����"O�����7F�6$��c^�nG�t["O��h�m�����Ղ:+�����"O�T����i��ȅX�	�F�q$"O(PS�PA�n`��23��|�`"O�w�/=����C ��[O��zF"O���d���{�I�D��5i��"Ox9��U)	�,�Q��!��3�"Ox�ha�Gj�����X��u"O���Q��큒�K�<s�x��"O���Q`IM�d�`��j�d³"O�"&P����s��=+�I3"O�Y� *[(�g�!��a�"OLR�dʮ0*����4M���"On�+�ύ=	��-��G�.2C���"O\�*W/F� ���<��"OE��ѹn�޵�r���^;*qP"OX��׮Ӥ`��3W�G,/+��"O^8qc��,k�M)U�!O*| qd"O\R�eQ\HpbR
�#D'F��"O�x[`M�p��䊳�T� �2���"O蠐B�Ԙ��Kw�V�V�v�y�`#D�`�e.E�-z�T�W��[CHI�+#D���GJv7�lZ�+��?~�}��C+D�d�D(C�{��(6!� ���>D� L�W����rE�M��y*��?D��ʲO�O��t���S=�-`uG<D��XUhͧTP,� s�?#-��v�&D���2"X�	�|0	��A'W亢	*D�tPg�ϨA���{4k 3��`���=D�@���<�v��g���!su9D�@qQ Å.0��w�
�pX�� �)D�$���Տ��� ��d�F�J��(D�8ke	کrظ��&Hd��8�e.2D����*F����j����@)�F1D��u�BIˑJ`����,D����`�/-eP@�(З�$lX +D�t���m����KA�< �&D�V�
�B�^�`�ϐl}
�Z�)D�,�g�?g�B���LHo����N;D�l�B�L�x�t,����*cc~hS�9D� B�Iĵp��es�D���%�Tn5D�� ���%�P�W�������>*?�� �"O���@npԄ���&!7����"O,�d�G�-��dڤ�ж}Ф���"OB����>�(,j��Ґ~�q "Oнq�!	5OXJl�tG
1[`z將"O~4�� *����R&��;Xb���"O`�a�Ǚ�Z�ؽ4_%l2��R0"ObP
$*ڽ7��Z��I�[��I"O�4��,W�z-lx�6��%$*��"O��KĎ͚+?~��[�)�q��"O�Iz&N�*̑E�\6Jٹs"O ����R7a�!K�h�!_
��x"O(�� �R�V�5ɟ�H^h��"O�(� lU%W�ʙ0�A��u���"OP���z����aəG����"O��.���ӂi�.6L�4"O�UJDW1��K�hݘQ�|�q"On�*D#�.�&�xdBرU` ��"O�Iz�e�?�h��!�~ֶ#�"O(]�$hR�wx`S��Y�'3��	5"O��Pl Mb3 ]�"�,��"O^l���ԡ	Wl�&n9L�[r"O4l۠�Ċlq@�u��$P-�	�"O�聄�#b���(�`X��̒�"O�����v'�A! -@ w"O�-a B�%'�j���G���G"O2;Df�b�\ذ���0ݣ�"O����Z�$���tN/�\�+c"O���`kA&��kʫ^�p��D"O��)AΚ�sX`D2 W� �D��"O.��g�>vAd�Z>&��Mhq"O�a���Lt]�ԥ'��ѣ�"OTъQ�R5KJ�((�dԷ@{�I�"O��S�LF�n�K��H�j ���"ObdB�MK��	�j�
gT��&"O�MhB'\�U�!�� S�4�H��"O���H�����g��g�
b�"O�ȇ#��$���
�0���"O����ҥ0ش�%��kVd��4"O��S
@.�f��ee�'\M3�"O�<(3Fog��8V%4,&�$"OV���?<z`I��ʶ{D{�"O֠���9v1��i�3`]�9�F"O���L*�L�X�)����J�"O9�`W�>��r�\��@q�"O�%6-zN���iU�� ��CVk�<ْ�"=����BC�j����% ]�<	��O:A]�L@d�M�!��qؤ��[�<)se�,jL���	TPjuG��U�<1�S�U�[rE��XԖcU,�Q�<��%�2�ճs
Y5i�B���TQ�<��]���*gmYbxP�[��y"
�oPL%�A#��Y
p�7�yB�Y�E%&X�ł�tl�Zd.U�yr�^�\;8Y�M7E�FE��y�:1N�-a�U(6j�l�4�I,�y��=mZ(��d��w0|tA�1�y�	�N���:{G������y2I�=�,���"r�D��tL�yB�D�2�:�`P�Þ<Τ�⭄��y⤅�m=l����boܰB��P��y""�ZDxR��~��ފ�ymƁc�IshP�9������y2-F(F�8հ&j��B�p��1�y
� HpA�P�=�N)�d �"�˄"OX�;�ǃ�D��b�̘�C��Xu"OȨ�&a\�w��RtƇ�*�zD�#"O�A���'x�Ԛ6eˌ�(�"O��P`E7Gb|C�j�-�
���"OԸ�$& ���n��l��"O�rWA�\f��O�'+�>�ɤ"OZ��Fo�.��n��e�dY"OL�����@�aS�ʝ�Zb��̺	phz fX�ęEE�
{�58e�ҩi��b+4D�\�V�R�^� ���P�K��ꖭ2D�Ti�=^�b��g==��y�2D�4��oa��z��K!�|<��.D�|�0�?p�,a(�%���rr�-D�Â*ߊ[�p��]�X���,D����԰,B�cE�:A�I1�,D��8�	;��e���/�/Ya�B�I%�F�i�MٮO�hЯ�K`|B��'J(��A�A�Cߠs�F�o�\B��#W5�y÷�NN0v-84�N[�JB�I�lDԑ��!����S���w�B�+�1��h���� ul3w�B�	�^=H!�c�p-��8תʰx��B�ɝ?q2��E����%��[*nC�I6;��<��,��ze�����D^��C��/*�!��Ʉ�U%�F��C�	O���c�NE9+q�f�Y�kA�B䉶xG��V�$�b�ؖ��n�,C䉻^�p���#1�F���a�H,C��K�v8!�@3 ]��[&��O,�B�	'xBNZ�N'O�9 �l��B�>���gbU$<ԐP�1≥4 �B䉶O0�h6�͑S�bP���u��B䉸B�z��%@L:�fѓ%�عgN(B�	�5�1r#%S1bf!2b��+JC�	Oy�pB���Ş�ӳ��cxC�	�-Ϡ�!�K�0]���	B�:��B䉃�]r�l��wq��B_=�C䉒ax@���.T�3���G�B䉖
Ք�� ș�7BԒ�@[�} B�ISP�)�`V,	],�Eb���C�ɹD���C��I5V�ءp�,��n��B��!k�hrum�S�Z4���Y8�B䉵fH�A�F#D�܄�5,�d��B�I�1v��� �Ĥ �kz�B䉾`�Ry�/
N��4���="�rB��e�
��FFͬv�丳`�>9�NB�I�� \�b�&�>��ƅ[ �B�I��J�[�`KV�6��3��~�:B�
^�d�Ѐ)�)M� �Ȝ�x�B�����ڄ-�(�$���Y�wB�I1k��h�)l��p#�
>}�$C�I-|�L�u/�PV���w�_��C�ɘ hxH���Y�`qL�AU	 iC�i�NA�tHmS��O�h��6�"D��+���?��$A#�
i>NTѢ�$D�@��
D37�f\dȐ\O���� D�X�%QG��٠�h*m�����<D�$z�(U�P.���� �6zr��Ч�<D�x#S��	8�l*�k�d����7D�X:&�ӓ%F���Q�Q�tppDO7D��I��L�BB$E���d��U	0�1D����D�TC�EQS�"g�Xq���0D��H˄�"�(tFC�R9���0�#D�� 
�aӭ���=��o��wb�S�"O^��\�f7����A�*��"O��ц �
��9���M q�6h�6"O����C�1��W۬0��I("O�j�jV��l�M]%J���ju"Oh�9�S]�`5�5,&���Bc"O�p�
U��P�C�'n��1�7"OԽ�J�f�21(����k��<��"O*����?3�U�Ţ_'XvĹ"O��ce�ڑr�Q�ա�:#u�;�"O�<��ca��MQf`�!Y���"Or�s�Fӿa�������#h�H-��"O
�2#��,&ޱ �D(�Jmj"OV��S�!P������g�i
!"O.0�ԅ�,I�(����D3���A""OR�Z��+�����ʃT�~]K�"OƑ��O.]�XV�̝^�ܣ�"O
4��i����ʙ43&Z!f"O�M{�F!Eh�3CoF� ��=	G"O��g�؍"�
\�Ү�d�0�ʧ"OZ	`��/F��A�SOI�3լ��q"O�ѻ`�NDZ9r�cF�c(���2"O ��7+�.K������9q$v	z"O"�Bӿ
�~9�F�N���[2"O6ə��(�|u�W�X�(�ّ4"O���tfϭҲAv,
#y
�S5"OaV�Q- ��쁍d�A[�"O�[5oN!\L]����!�;1"O�b����a�R�A��\��$y�"O�C�i['e�p���h�7�DK�"OTTS�Ĩn��AP�� )�|AP"O�� ���jӎU��/d��8"O0�)�A5����wD��ey�|Z#"O�%r4�V�
�����I(D��\��"O�5��F>�����C#n�RЋb"O�qi���$?N�A� 5���C"O����-vrɲ׊I�,���"O���Ԫ�|,8�:��ȫ{
]q!"O ��:"�mc��N/Ac-"O>�Z�,	*R� �G(O�Pb��RA"O��!�b�X��g��|+���"O��s�"1�@� ��L�U�v"O�͢�j���\B���<�)��"O<����B!\�<aQI�(|�P�"Oཱི�N�]8�(��$b$"O虘%!�!UX�=�㇈�T��ZR"O�4z��N+mEB���睕 Tu��"O�� � ��dr��	~׸Mr"O�TQb@�M��)+��3"��T"O��;B/�]��iYĎHl��@�"O�a��&W-S$>M	V�><j�
T"OH��E	�/)ˀ� �
K8<#�P"O�	p"IDq��P���O�7q�i2�"OX�æƪ:���Bi3N�L���"O��d ����V��f�A��"OLX�b�fbLPIU�S�D��"O�%��Ǘ*�TPHϜRd@*�"O���&-��8LƝ7�¡aF��P"Ot0k7PE^h���ʎ�jM�"O�q�E
�#5��j��}۲a:u"O|��+$-����/��P��"O�I�ǠM�L�&-�"Q����'"O�A�`�ִ\��qo�e���{�"O6�#`ʋ>N &�eo���Ac"O� v��B�8r�m8V���>L8 �"O<t�sŃ'W��Q��r=��9"O��z�I�/!		(�̇+
1
9��"Oū"��GB��'뚡B$*��t"O��4��G��p�i��2�AT"O��E�S�:8
C	��P��"O��:c�>W�Q4H�$�L�d"O6������Dk!���̬ct"O��P��ce�C	KR4���@���y�M�/D~�	v$
�B����G�C-�y2���(�Z��������yB/A�! ��D/Xw�>���H���ybD�x@��P���z2�$�!.���y�CV����cx�F�A��y2�Ӣ;���f�}ü�� J��yr�4~�b0IdGL
,|8��T��y�͒3f$�я�Sz��Ў���yR���rbN�:UdҢE��i H���yR�åu���TD�.A2��F�<�Q	�<�0��5*ؗs��9�t�<�@��"�����k�>���e�<��FU���𫘅F8`�SX�<����&c|�A��F)޴�����z�<y�, $����_#c�E�2jQv�<��A�. �d�H��ߕ"=l���q�<�Ğ�+��9ro*	z�u�Bʃp�<q�_YP�0xf&�X�(�T�<�%i��<���r���1�}�A�R�<��-P����c�-O�,���c�<���ϘA=�p�4O�_R,���C�<�ь�9\%;��'Oi�q���C�<	RI�p�TYCq����Z���t�<qO )���`ԍ=^��R�f�|�<�c� 
�.t��Ɔ�������z�<��F�0`i��;��^���ȥ�x�<a��ֺ55Ό��>a�Qx�ΐr�<i�Ɨ,"I�˾$�AXr�Hi�<��iI�6P#׷)�� �#�y� 2P �	7@šqg�<��K'�y���K
̻e�?a�cA� �y�M8��#�YF�P[a �;�y�晃3��"s�#$��<�͈=�yb�R̢��i��^�c���yrK�(�$8B�
�ެp7ƅ)�y��ſ7�h� ��5�Yk���0�y"�Z4<�(c�јx���xФ��y¥�������ݕk���	����y�V%d��A�A]fhɥ儈�y2g�6|c��#6b
�~��S�y��6��H��._�ze���@�P��y�.�=����l��QkE�y�υX�\(w�`"�j� �y�M� \�<��CU)`�M	�y�AY#p,<��b��?R��A ��y�`S p�c��*MJ��[�N��y�Ӈ$Tx���5Kb������y�nZ*	�t����:2�I�F�G�y���~ ��ͻ+n���fF�yҀ ,A�D�#'iI)s�F�!׬�y2�YD�ɠ� �=��8�M�)%!�D�a��H��� �aZe�G�!�-IDQj$U���@�ƽ/�!�d[4IT�p��<G���a�*)&!�َz�h�E�ӊ3Y4�J��ly�	��� uJ�e��@9(H �j�&�|��"O�H�W#U����ʄJ_�����"O����)){��Q1G��|x�m��"O��)R��K
̨䥛:;u±q0"O�����ވL� �W�VV��Xu"O�0��/M�`��E�&�.�%"ON���M�\�BɻvB6A��@"Of�J�^(d���PJ�p����"O���.I�LqK'���o�� ��"OȄHP� �	X[2�p٣G6�ybgH&Ŧ	ʄ�ь{<�##Ώ��y��W<US8t�C�y�����ݯ�y��Z�pg��% P���D�>�yR��~   �   6   �L#�靱I����t�B��L�:�.ħ�~��'(R� e'�(���(H#b��!�o�|�d\�+�yK0l��~����c��83F��m�5�M�%�i�r��$���H���5K���'N�����቉U���3A�i*�)�
B�sBD�ai�68dEr(O�q�TI��<@��`UX��{D@Z,�� �´>!���85�fT���y�J�9�T�\�If��m���<v�@�WF�}���9lB�Hh�@J�b킧o��r:�8�!���F�4�ɠ|�?Op��
E�:>r�y��{L�Z��|Bc�'0�&�D��k��0Q�욅��HZ��'�}�4
��	�F���@��7`�F|�ާs��� !a���OڭI��d[;��D��[; ���,��}ź8����)F��t"<qV� �	;��V�S�9j� #��
�j6�\��Oޑ��d»�H|0�A�>
�Q�5a*�2��$X�OV��O$e���P��,�c���F�r�1RP����	4��O��臭�E��"�+n�2	C��O�:���ӂ�?�w㋊m����� _���*&͇p̓ �"<��%�I,zRi��&�]�PZ X����O��8�y2�	�kz*d+w��L匭� �W�5,0��r�'v�(Ʉag��pʏ�Q����>���&2�Ш�	ai*1PB�/4�؀5`�&t��t��ɇ.��.o�����A�/�z�QrB9uo.M�'�Fx�i�'s���4fy#��p����'ePPY@ ��lh" M�6�6@�%?:��D"P���V��R�$9e�.)T$�V
O���ֆ`ӾLm<60�'�@�`,z�r%ɓ�0#�FCpdPq��i�R����Gڟ\��&��d��Uܣ�~��BfCԟ��?)B�Z91�fe� ��T�X�	B/h��Swi�b!���j�vin��?	�S��֘�"��3��8;/va��ވl'2���ۘTT�}�ȓ~ȴ�C�O�H��*g��g�jцȓ=�vL+��'B"�HHf�]�FB��//����N:��`�

eG"��ȓl�j�ړi�`1��H���
���{��-3���0uʸ}�Q��<NqMD{�.�����l$�D(�b[����
�@�pa��"O4p��&�7z`y��1$��=�4"O�7�."t0@f��<3�0Rd"O4�5!ً2x!�,�?i�&"O��¤�2:\u;�    �    T  �  �  '&  y'   �L#�靱I�8��tE*���"O�$��L�'bj�����΂<4��ش"O�Ȩ6���U8�	���*�)���o�� #��4h0�`Ü�b�ְP6�	;D֑#�����g� s��q��,I�A��Q*��;d�����g�z�g��D�tq��\�WOB��&)B�m�1���/L���4��{���93�N#7�e����~Y�A�(ۚ�賠�YX����*�$�N����,\��0��M&D�����, n�e���R���0Rqc0D��i��J2?�e���*���u�?D��e�Ӥ9HJ$���X��dbL"D���A�(s�ZvKP.�H`H!D�������z@��34̀S���p�#D��a�'[�8`�v�D�*�q�4D�����8O(�ҒOU�ra�0ѷj4D���5���F����%��!i���m1D��8t�M�rJ|����"c���)D��n��'ep`�W�S~(����6D�PZU�]Qg8-�j�#/N�d�5D��`�	֋q3�����n��4D��ڀ�S.��ԁi�)�ZD��7D�LⳄ�
�1��L��<�d��#D�hr��)_ �5!�''Ҡ)�g"D� 8�Ʌg�1���-G���xeN%D�<�`Q�91����+����b"D�@��;^s$�[Ѝ�24���d�<�գA�%c
`A��B
L���0��C�<`���J�S�)@��̩B��g�<���&'�n(dj��H�h�M_`�<���{�#�W�e���s�`�<!�g�BG��R�,�<Fjl�Y@�y�<!l�=k�R��#�=)�@��%�v�<���I'PѾ��F��/W�4q�E�s�<	A�	~�&xQ�	�Lr 9qQj�<�VJ�֭���$��XA"Cd�<���;Q@�1���E��d:�i�<�B��Pa��3�$2dt$�N�<�gg�
�L�!�	�0BԄ�A�@�<���U&�ԭ��mX
 #*���"\v�<a��7ۼ�蓫?U�(,�@ v�<���U�|�H��#j���SC�Pr�<v�*lj�+u�H0�Ri�X�<Y��94���1� �r8�"J�<���ʋq*t���4<�`�Y�"�E�<i�NB�Cy���5
�w�r .C�<)5�>q��S�c̙�m���D[�<�Q&�/ ��YD��<^P��siY�<�ӣ�`fH��FcU9EP�+�S�<a�Ԋ�Dѳ�E�z��)q'{�<����!eƮف��݂W%x����m�<��ʓ({�nPD ���T�`�<��M5�DȒ� z^��SE��<�4�ͽ^U�H ���<��]�5�Cz�<�w��i;i�ɟ>5�23�"	s�<Y���.D��3A��8����N�O�<d�أJ�(b���i���A��YM�<Q�H^Myޱ2�bZ	%B�32��O�<���%m�r�2���/b:Ղ���p�<�gύ�<�Nq2��O�L)��B�M�M�<u��V��M��`ˊ;_��0A@�b�<i�B�pb�MA(��4)H|��EX�<��MW��p2���y��U�<�#�+9��� $ڋ5N��F&{�<Q%�U�?@V#J�A�H�jD��u�<a�fR1]�L�QN�QJ-���y�<�lG�=	��r�lV�f��BOPx�<� ���Ec�b�pyy�m׍J�����"O�@�V@ό#+���"�WG���"O�T�`�ۊ�Jp�p-I_�����"O(�A��:��	q�R'K(��"O�M:˙�d���Bu����"O^��l� %N5	"�m��(��"O Y�B�E##��r ���R~ԁC�"O��G�Z�.�^�����8Met0�"O�Yy`E>J-��d'F(�"O4�B��B��ݻ��W�1���Zv"O�,���K,o��ٸ�I��h�,�3v"O�$I�krQ�"*�K6��"O�j��B�L�����;7"H�[�"O ��X~C�鉷��'f��!�"O��
�b��=(��\�C&"O(���c�\�5��I�'J��4"O��q&b,�Ŋ��^���R"Of%bY5�v��6%��e���`"O|���ف+����a��3�`4��"O(� ���)/�a� 3�����"O����ѹ0���⧞�n��d��"Ot=㱪�t���+� E�*vmش"O���g	�;{�0���G�*Wb����"O�����7F�6$��c^�nG�t["O��h�m�����Ղ:+�����"O�T����i��ȅX�	�F�q$"O(PS�PA�n`��23��|�`"O�w�/=����C ��[O��zF"O���d���{�I�D��5i��"Ox9��U)	�,�Q��!��3�"Ox�ha�Gj�����X��u"O���Q��큒�K�<s�x��"O���Q`IM�d�`��j�d³"O�"&P����s��=+�I3"O�Y� *[(�g�!��a�"OLR�dʮ0*����4M���"On�+�ύ=	��-��G�.2C���"O\�*W/F� ���<��"OE��ѹn�޵�r���^;*qP"OX��׮Ӥ`��3W�G,/+��"O^8qc��,k�M)U�!O*| qd"O\R�eQ\HpbR
�#D'F��"O�x[`M�p��䊳�T� �2���"O蠐B�Ԙ��Kw�V�V�v�y�`#D�`�e.E�-z�T�W��[CHI�+#D���GJv7�lZ�+��?~�}��C+D�d�D(C�{��(6!� ���>D� L�W����rE�M��y*��?D��ʲO�O��t���S=�-`uG<D��XUhͧTP,� s�?#-��v�&D���2"X�	�|0	��A'W亢	*D�tPg�ϨA���{4k 3��`���=D�@���<�v��g���!su9D�@qQ Å.0��w�
�pX�� �)D�$���Տ��� ��d�F�J��(D�8ke	کrظ��&Hd��8�e.2D����*F����j����@)�F1D��u�BIˑJ`����,D����`�/-eP@�(З�$lX +D�t���m����KA�< �&D�V�
�B�^�`�ϐl}
�Z�)D�,�g�?g�B���LHo����N;D�l�B�L�x�t,����*cc~hS�9D� B�Iĵp��es�D���%�Tn5D�� ���%�P�W�������>*?�� �"O���@npԄ���&!7����"O,�d�G�-��dڤ�ж}Ф���"OB����>�(,j��Ґ~�q "Oнq�!	5OXJl�tG
1[`z將"O~4�� *����R&��;Xb���"O`�a�Ǚ�Z�ؽ4_%l2��R0"ObP
$*ڽ7��Z��I�[��I"O�4��,W�z-lx�6��%$*��"O��KĎ͚+?~��[�)�q��"O�Iz&N�*̑E�\6Jٹs"O ����R7a�!K�h�!_
��x"O(�� �R�V�5ɟ�H^h��"O�(� lU%W�ʙ0�A��u���"OP���z����aəG����"O��.���ӂi�.6L�4"O�UJDW1��K�hݘQ�|�q"On�*D#�.�&�xdBرU` ��"O�Iz�e�?�h��!�~ֶ#�"O(]�$hR�wx`S��Y�'3��	5"O��Pl Mb3 ]�"�,��"O^l���ԡ	Wl�&n9L�[r"O4l۠�Ċlq@�u��$P-�	�"O�聄�#b���(�`X��̒�"O�����v'�A! -@ w"O�-a B�%'�j���G���G"O2;Df�b�\ذ���0ݣ�"O����Z�$���tN/�\�+c"O���`kA&��kʫ^�p��D"O��)AΚ�sX`D2 W� �D��"O.��g�>vAd�Z>&��Mhq"O�a���Lt]�ԥ'��ѣ�"OTъQ�R5KJ�((�dԷ@{�I�"O��S�LF�n�K��H�j ���"ObdB�MK��	�j�
gT��&"O�MhB'\�U�!�� S�4�H��"O���H�����g��g�
b�"O�ȇ#��$���
�0���"O����ҥ0ش�%��kVd��4"O��S
@.�f��ee�'\M3�"O�<(3Fog��8V%4,&�$"OV���?<z`I��ʶ{D{�"O֠���9v1��i�3`]�9�F"O���L*�L�X�)����J�"O9�`W�>��r�\��@q�"O�%6-zN���iU�� ��CVk�<ْ�"=����BC�j����% ]�<	��O:A]�L@d�M�!��qؤ��[�<)se�,jL���	TPjuG��U�<1�S�U�[rE��XԖcU,�Q�<��%�2�ճs
Y5i�B���TQ�<��]���*gmYbxP�[��y"
�oPL%�A#��Y
p�7�yB�Y�E%&X�ł�tl�Zd.U�yr�^�\;8Y�M7E�FE��y�:1N�-a�U(6j�l�4�I,�y��=mZ(��d��w0|tA�1�y�	�N���:{G������y2I�=�,���"r�D��tL�yB�D�2�:�`P�Þ<Τ�⭄��y⤅�m=l����boܰB��P��y""�ZDxR��~��ފ�ymƁc�IshP�9������y2-F(F�8հ&j��B�p��1�y
� HpA�P�=�N)�d �"�˄"OX�;�ǃ�D��b�̘�C��Xu"OȨ�&a\�w��RtƇ�*�zD�#"O�A���'x�Ԛ6eˌ�(�"O��P`E7Gb|C�j�-�
���"OԸ�$& ���n��l��"O�rWA�\f��O�'+�>�ɤ"OZ��Fo�.��n��e�dY"OL�����@�aS�ʝ�Zb��̺	phz fX�ęEE�
{�58e�ҩi��b+4D�\�V�R�^� ���P�K��ꖭ2D�Ti�=^�b��g==��y�2D�4��oa��z��K!�|<��.D�|�0�?p�,a(�%���rr�-D�Â*ߊ[�p��]�X���,D����԰,B�cE�:A�I1�,D��8�	;��e���/�/Ya�B�I%�F�i�MٮO�hЯ�K`|B��'J(��A�A�Cߠs�F�o�\B��#W5�y÷�NN0v-84�N[�JB�I�lDԑ��!����S���w�B�+�1��h���� ul3w�B�	�^=H!�c�p-��8תʰx��B�ɝ?q2��E����%��[*nC�I6;��<��,��ze�����D^��C��/*�!��Ʉ�U%�F��C�	O���c�NE9+q�f�Y�kA�B䉶xG��V�$�b�ؖ��n�,C䉻^�p���#1�F���a�H,C��K�v8!�@3 ]��[&��O,�B�	'xBNZ�N'O�9 �l��B�>���gbU$<ԐP�1≥4 �B䉶O0�h6�͑S�bP���u��B䉸B�z��%@L:�fѓ%�عgN(B�	�5�1r#%S1bf!2b��+JC�	Oy�pB���Ş�ӳ��cxC�	�-Ϡ�!�K�0]���	B�:��B䉃�]r�l��wq��B_=�C䉒ax@���.T�3���G�B䉖
Ք�� ș�7BԒ�@[�} B�ISP�)�`V,	],�Eb���C�ɹD���C��I5V�ءp�,��n��B��!k�hrum�S�Z4���Y8�B䉵fH�A�F#D�܄�5,�d��B�I�1v��� �Ĥ �kz�B䉾`�Ry�/
N��4���="�rB��e�
��FFͬv�丳`�>9�NB�I�� \�b�&�>��ƅ[ �B�I��J�[�`KV�6��3��~�:B�
^�d�Ѐ)�)M� �Ȝ�x�B�����ڄ-�(�$���Y�wB�I1k��h�)l��p#�
>}�$C�I-|�L�u/�PV���w�_��C�ɘ hxH���Y�`qL�AU	 iC�i�NA�tHmS��O�h��6�"D��+���?��$A#�
i>NTѢ�$D�@��
D37�f\dȐ\O���� D�X�%QG��٠�h*m�����<D�$z�(U�P.���� �6zr��Ч�<D�x#S��	8�l*�k�d����7D�X:&�ӓ%F���Q�Q�tppDO7D��I��L�BB$E���d��U	0�1D����D�TC�EQS�"g�Xq���0D��H˄�"�(tFC�R9���0�#D�� 
�aӭ���=��o��wb�S�"O^��\�f7����A�*��"O��ц �
��9���M q�6h�6"O����C�1��W۬0��I("O�j�jV��l�M]%J���ju"Oh�9�S]�`5�5,&���Bc"O�p�
U��P�C�'n��1�7"OԽ�J�f�21(����k��<��"O*����?3�U�Ţ_'XvĹ"O��ce�ڑr�Q�ա�:#u�;�"O�<��ca��MQf`�!Y���"Or�s�Fӿa�������#h�H-��"O
�2#��,&ޱ �D(�Jmj"OV��S�!P������g�i
!"O.0�ԅ�,I�(����D3���A""OR�Z��+�����ʃT�~]K�"OƑ��O.]�XV�̝^�ܣ�"O
4��i����ʙ43&Z!f"O�M{�F!Eh�3CoF� ��=	G"O��g�؍"�
\�Ү�d�0�ʧ"OZ	`��/F��A�SOI�3լ��q"O�ѻ`�NDZ9r�cF�c(���2"O ��7+�.K������9q$v	z"O"�Bӿ
�~9�F�N���[2"O6ə��(�|u�W�X�(�ّ4"O���tfϭҲAv,
#y
�S5"OaV�Q- ��쁍d�A[�"O�[5oN!\L]����!�;1"O�b����a�R�A��\��$y�"O�C�i['e�p���h�7�DK�"OTTS�Ĩn��AP�� )�|AP"O�� ���jӎU��/d��8"O0�)�A5����wD��ey�|Z#"O�%r4�V�
�����I(D��\��"O�5��F>�����C#n�RЋb"O�qi���$?N�A� 5���C"O����-vrɲ׊I�,���"O���Ԫ�|,8�:��ȫ{
]q!"O ��:"�mc��N/Ac-"O>�Z�,	*R� �G(O�Pb��RA"O��!�b�X��g��|+���"O��s�"1�@� ��L�U�v"O�͢�j���\B���<�)��"O<����B!\�<aQI�(|�P�"Oཱི�N�]8�(��$b$"O虘%!�!UX�=�㇈�T��ZR"O�4z��N+mEB���睕 Tu��"O�� � ��dr��	~׸Mr"O�TQb@�M��)+��3"��T"O��;B/�]��iYĎHl��@�"O�a��&W-S$>M	V�><j�
T"OH��E	�/)ˀ� �
K8<#�P"O�	p"IDq��P���O�7q�i2�"OX�æƪ:���Bi3N�L���"O��d ����V��f�A��"OLX�b�fbLPIU�S�D��"O�%��Ǘ*�TPHϜRd@*�"O���&-��8LƝ7�¡aF��P"Ot0k7PE^h���ʎ�jM�"O�q�E
�#5��j��}۲a:u"O|��+$-����/��P��"O�I�ǠM�L�&-�"Q����'"O�A�`�ִ\��qo�e���{�"O6�#`ʋ>N &�eo���Ac"O� v��B�8r�m8V���>L8 �"O<t�sŃ'W��Q��r=��9"O��z�I�/!		(�̇+
1
9��"Oū"��GB��'뚡B$*��t"O��4��G��p�i��2�AT"O��E�S�:8
C	��P��"O��:c�>W�Q4H�$�L�d"O6������Dk!���̬ct"O��P��ce�C	KR4���@���y�M�/D~�	v$
�B����G�C-�y2���(�Z��������yB/A�! ��D/Xw�>���H���ybD�x@��P���z2�$�!.���y�CV����cx�F�A��y2�Ӣ;���f�}ü�� J��yr�4~�b0IdGL
,|8��T��y�͒3f$�я�Sz��Ў���yR���rbN�:UdҢE��i H���yR�åu���TD�.A2��F�<�Q	�<�0��5*ؗs��9�t�<�@��"�����k�>���e�<��FU���𫘅F8`�SX�<����&c|�A��F)޴�����z�<y�, $����_#c�E�2jQv�<��A�. �d�H��ߕ"=l���q�<�Ğ�+��9ro*	z�u�Bʃp�<q�_YP�0xf&�X�(�T�<�%i��<���r���1�}�A�R�<��-P����c�-O�,���c�<���ϘA=�p�4O�_R,���C�<�ь�9\%;��'Oi�q���C�<	RI�p�TYCq����Z���t�<qO )���`ԍ=^��R�f�|�<�c� 
�.t��Ɔ�������z�<��F�0`i��;��^���ȥ�x�<a��ֺ55Ό��>a�Qx�ΐr�<i�Ɨ,"I�˾$�AXr�Hi�<��iI�6P#׷)�� �#�y� 2P �	7@šqg�<��K'�y���K
̻e�?a�cA� �y�M8��#�YF�P[a �;�y�晃3��"s�#$��<�͈=�yb�R̢��i��^�c���yrK�(�$8B�
�ެp7ƅ)�y��ſ7�h� ��5�Yk���0�y"�Z4<�(c�јx���xФ��y¥�������ݕk���	����y�V%d��A�A]fhɥ儈�y2g�6|c��#6b
�~��S�y��6��H��._�ze���@�P��y�.�=����l��QkE�y�υX�\(w�`"�j� �y�M� \�<��CU)`�M	�y�AY#p,<��b��?R��A ��y�`S p�c��*MJ��[�N��y�Ӈ$Tx���5Kb������y�nZ*	�t����:2�I�F�G�y���~ ��ͻ+n���fF�yҀ ,A�D�#'iI)s�F�!׬�y2�YD�ɠ� �=��8�M�)%!�D�a��H��� �aZe�G�!�-IDQj$U���@�ƽ/�!�d[4IT�p��<G���a�*)&!�َz�h�E�ӊ3Y4�J��ly�	��� uJ�e��@9(H �j�&�|��"O�H�W#U����ʄJ_�����"O����)){��Q1G��|x�m��"O��)R��K
̨䥛:;u±q0"O�����ވL� �W�VV��Xu"O�0��/M�`��E�&�.�%"ON���M�\�BɻvB6A��@"Of�J�^(d���PJ�p����"O���.I�LqK'���o�� ��"OȄHP� �	X[2�p٣G6�ybgH&Ŧ	ʄ�ь{<�##Ώ��y��W<US8t�C�y�����ݯ�y��Z�pg��% P���D�>�yR��~   �   N   �L#�靱I���d�C= �L�:�.ħ�~��ק(R� e'�(�����G"d����l�<�dӿBRT��3c�/�f��v�S�TD�o��M˲�i1f��$�<(HQF-( �ǂ0����ቝQ����õi-x��م,*6�H� �5���+On`��G�84�#]�P�A�|��욂oo��!-���(�
�N�4p@��B�5A��EP�rٛ��O�扞"�<jҽ�=b-O�ԨB�y���d0�64h��;4���-���G�_}����DPx��II���)F��5�kW0��e��!Er�H`Bא1���$�xK��1o��'L2 3J�>)1huj� �90&��H�'\�Dx�KA�'�>Q"K�t�T=xᤞ�b�����$MP#<ѵ�>��
�,�2!��f�5��*B�����O��ˈ{�lI�n�4A��)��nF�5�P�]�Ms��+�Z.D"<�A+�Z���P6�b�Ĺ2T�ە)���>	q�5�U!P�\���2­\�"��r/	'N�vM�'��@Ex�A�n��C_F8i�*eoؕ(`�W�V�X��;4x@#<Q���O�q�f;qr0�jv`��w�pA����O��O<�W*׈H[�pg+�>,�+��o?!g$�7�c� ɇ��~��e'#���¤��2.���`���:WG�9PJp�CF��M�J�0Ʉ�L������ZA6u�&.��v�@zUM�@<qO޼R��$���7obQ	U*Nn%d�&]!�:�-qT#<��1�<�f��0k2[�`ZGh���0�ȓ���  @�?�bDk�"��9��B䉇MF�PpԋD 4�&�"�a�TY�B�ɜ_�8��拀J�|s���F�B�N7��@��#:w�ق�&�vB�I	(����䑣��U����2h`B�ɚMxh�a�.'���	u�!} XB�	4|E��Ԇ ����K�(B�I2qrP�é�:e�A��-�2=/�C䉰hM,��1�P��H0jU����C䉫!Y��џ_���Є�>aXZC�ɳv�D��~���y��I�C�	�7���ۀ�T�P��bձ
ŜB�I�����&�DYH�E�8B�	(���1Q�4D��3��6HfB�		x��̊���2aof�r��e�XB�Ɇn�Z�c��\��qj��rB� i�(�C��1�N8U��!zC�	�Z �Ҡ�O� ,&�y�hG�B�I4c���'I�p#���r� B�	�xYAj7`@�oޜ 4�Bu�B�	"(�	��2
�f����>��C�	�Pa$���.��I� |���%�tC�t�\a0�ۭ8+҅��*'8�@C�	N�8��훡j�e�%_�D$C��
~�$EY5�_�)�ֈ1$��b8C�I-$��y{��A���8��Ghe�B��?;�R�s�.�=a�� *��J��B�I+7��z#��* ���iw�ǫ�rC�	�f�|��"!؜p&VL�@�C�lC�	,x��k�]�k�V��fB  ofC��6+i(r2i�[�X"Q���2�B�I*0�{�e��!E�����(&lB�	b�k��E�,󶴀��W�@S"B�)� ���2+M�v��s\�)X��T"O~�U�Ё��<���^���:1"OF����Q$�����'htD��"O�-�t$H��Y��kB�J���"O��!��?^̀EؠL�A>�V"Ov��D.X�t��T�i�.8��"O*��P"JBp�̂��P�}'$�B�"OxM�uM�&r��M��Ɋ4���"O�9�V�+$�ӳ��-n2L��"O����Y�p�T��"��c"O�Q�pƒSw\�3E�6�X`�'"O$m����%*R�hR�ބ���"O�}3"G7� 1�Ab��Dk�"O\�8P�G>��t1t ������3"O��ؠ�݊IJ}
P@]�U� չ�"O�j`��3Lڄ9t��8�L�)�"On��N��z���v��3��y�"Ov�� g��*����s�@D��u"O4��#�̷V,p4�Q�.\G(�#�"O`�(�`@�LJ�����.:�<��"O�myk�p?�Z���v�!�$7:Ƹ��	�>N r���D�>\�!�$0z߼�8������S��OPf!�䊪
l9�b�XC��Zq�_P!���?�*�c�̀�'�\RH�6Z!��
�D�+��� �>��Ԥӽ@Y!�&Y}��s�	j|z!5-ML!��@3a2�x���AþI��YD!�dO�|$B�ҤH�f�����Ǚv,!�$ԫT�u�P&7V�"��hأ1*!�d�o�u���H
ab�f!�d'��I�$��.�-ٶ�0!�X�<��mU-��B��vT!�;$V���S��R�h�ra׮cM!�$P�kV~���.(vc
53!�]!�!�䎊s���Sdc�5dGX��#o�T�!��'g�ذA�/6+�!�S�5a�!��\)-y^%��'C.�1NU�}K!�B�( ~� �N]&�m���ʷVJ!��˜��LX�X#�������?H!�§ۀ����vW�	�eD!�Ca�`A2A�<�ؽ�aOC?B!���&
m��i�o��"���qM�6�!�$�E�,���-�^���K�2�!����5���'������l�!��NcL�����:ݙ��V?e�!� �b��h�φ��t�Bだ�!��:8���9a�[7SQb��K6(!!�dV�:G�H����g��;�
[E�!�� �3��]��}�V�����8�!�䛭*gVH  Ѱ'4d$P4f�p�!��q�:1�7n�dƠPc�P=!���?��F�_*E�,�W�D�9@!�$� ��y�҆�pʺ8:���r1!�d�P� ��D�+���b���#n!�D�9����N��'�ڨ��D
<!�Dà_��:���5P��������!�Ě `���rE�J�A���BEoB]�!�D�p*�TxsϚ�H�� C�� �!��	�b�p�b��/(�hcw��30�!�d�?�.| �C%2f4z�oߪau!�D�<�rS&�Z�z��A$��d;!�..ZlZ ��w�jk�#μ&�!��M�f����g86ZY��� +�!�� ���˛�y���ce��%2p6�ؖ"O�ca�4?�hz�Y [v�1D"OD)"��I>�g��
gLM�t"Ox1��J�}�D��D�080�q�"O<�:B��L��E�̍£"O 8s���o��!��4���"O�m��P��`��D�9�uP"O�P�*�s���PD#�n�vY�"OM@v��=��-��a	)	�LPR�"O�@y�ړA�V(��T�L�ɓ�"On�Ҥ�X,��k�R���Y"O�	�Ǒ� T��KX"<���H�"Ox�i7b	qu�)� @��j��в�"O��1� I�Y^683�&Q�T	��"O�1��M=�#�/�8S
�PW"O$����"I�$�է��u��Iy�"O����Q6re�w�^�	�B"O����g�!|=:p�`Ű9!q�"O|M�d�!�^���;a�0��"O8M�d�?o�TUQT��^�y�"O�8��`�*�$8�7��2O�0���"OZ����+<;�ϓ�A�<�q�"OHX)�Γ�|x�C�N5Q윹"O��R�֙E �h��,�F�L�"OR�F	J�J���G��0QC0`�"ODZG)�k��I����C&�XP "O��)�S�:�T���G �as�qk7"O�5��.�8�D��t C�1\��8�"O��1��y�� �$n=��b�"OԵ��%��s�E�:
/���4"O�M;��pN�9`N�r��qyR"O���$Ҹ<�97��.ܘ�9f"OhY���9	hL��L��S���`"Oց�����X0��Ĩ�A�,I�&"O4 EÍ�lbL�;R	\�Xd'"Of�wHC�d��|��hT��:]�g"Oؐ)�� ʆij�7j��)'"O�%��!�%_��`$=(8A�"O��g(�	IA�i	�kY2G� �"Op\၁�*z�7��ns��b1"Oh��%� 1�(pɓiК`n΄1b"O�e �FI+9N�;��C�k�ru"OH������\�l�p���!/(�"ON�jP��Q"D���V+h 0�"O<�zR,��1\t51 "O��c`.�W6X� KҞ����"O�D �D�-O�Y��	�p�l	2"ON��S�P�W�V@9�i�?��PS"O���� �o��s���s��AK�"O�2�XwvT��� r��2"O&� �&�N�}��)Y�Y<"���"O�)c
��e���Ã܄.3)� "O�(3 ��Y��5�H&��h��"O�T��U"j����Ä]��"OT,A�O��?,h2� ��T��"OZ}���]�t���I��N�p�i�"O�tI�@Ap��yR/��L�\8����G�Xn��5�C
$J���6ɛ�X�'�N�A㖔n�*Ȃ�	�4L�-�
�'$(%��c�X�G��J�µ*
�'�
W"�(/X�$�6��BN9	�'�n5IUL�]�ސ�VN�6�-��'�ry�e�{�fM���6u{`Ab�'�們m�4���a�>^�F�!D��;��ģF�8���CA��Qa��4D�� *�Є [	142aBᦊ2[��	SP"O��Җ�[!5β�*��.+��4�"O�h�&��6�x�XbJ�� �*���"O ��E�!�������0�\��"O��ADB�k����!�Ii޲*Q"OP��e� K"^`�7�q��훑"O��ҧB�E�Aa6�]���lRQ"Ov��LB�u�H}���XeזLZ�"O��у×�O�X��-͛R׀�c�"O$��	��h;5Mل̠Y�"OJ98�E�6�0m��f<)�#�"O��%��z�:l����G�АT"Ob%��c��\��騠i	�˦|�D"O�(�'��?D����O�J:Ƶ��"O�3R�L(u�v���.�5G~�a"Oԁ��eg^!��Y��j��A"O�0D��6B^``�3ˑ0z���"O�����U7İiX����M%� ��"OJ�zuIH�d�x�u%ΫVN�b"O�8�I),�t�"���O���s"O��X$�:P`�i�td�	.�`�"O��֪��,�0H����q$�J"O�e;&d��:��P��l)6 2�)E"O�1��G�����N~5����"O"y�U(6k��Ԍ
eL�� "O6����9q4ɚv�	<���q""O��1CԸ}-�����'p��"O0���͋��r��e��wa0p�A"O���f��*F����%v-��J�"OD����ߥ�B�	�$��m��\��"O��v��.Ih�=�g%�Y~���"O]�IE�&H2ċ[�of�}ѥ"O����ڬh���S�+��>_�� �'|����?F 
�ȟ8'P�q��'V��F��*t`n �uN�uT��'�<5j4D�9t>�J�~���I�'����H�
μ [sJ�&��	�'.��& ȍ+����ϑ�"NJ��'!:D�O��\��0�Ah���'�[��V�1�8rD04P��
�'�N%*U��}���HE�T)v~�?D��'�q�HB�	Z�y�5D�<����1�n�BWG��Ir�2D���B�����{B�Y"\���a0D���d�و:�V\�!Q^W(�Y�F,D����օ '�xF�J ,.���C+D�tj�L�z�jI@AN��V����7D��;�&�b��ģ�I��X�x��A#D�,0 �	��y��	�7jBT !D�4�&L�}�(쫔�	�"�fhy!B!D��c2� @f'M&B P�� D�pz��z�f�1@�͋p�����0D� �Fb�8&@eaӇ�Ix����=D�(Db��?ZT��`o�i:��Ӆo=D��9D#{ �Q�ݲJ[�$�V'D�
���i����O�&pjii#c/D����]�"3�K)	���`7/D��3a�*l$p�$@W1!.@,bW� D�����C F�0�3Ƒ���p�c@/D�p{#
�Z��Aʑ�̀Q�n�`�,D�h�dLJ$����C˅5���'*O����K3�i����9@�"O(:����z:2#W�S���@"O��*a�
6g�|(��o�\��q"O�  a�"�)|<R���"6V	��"O"��@o�x(��B�~M�t�"Oք�b�Ĥ[�l4���E�]��q�"O��E�җW�P�锎�>,�>���"O���]�c��U�W�]�i�X�pW"O AZ�Y)>�I�lٜ!�4�"O�i��.L�qTu����Uq�"O��kV Q���k"<��,��"O�%�	5l�%H�,�-N�H�[�"O��1֪C?lR�h��Ι)���D"O��[b�V$:��á������G"OP�87�]0�0��y��	+��(D�����D�K�X7o�]�7�2D�p�S�+�ؙA���#Sh|�+D��NK2z���mЩ�&y걮*D��CrB�b��Ph&�ݫV�	�r(D�p`G���1��O[ۊՙ�6D��5%��x�LT��'1�� ��3D��� ƫo�H����F�>\���I0D�T�uC�E�4yG �0%��A�l?D�pG
P�z`U-^�Q�n���(D�����g�| ��u�۳�7D��A�O�94j�$C�_�<�e32�3D�Hr "E/�$0$��Xt�IR�0D�"W�I;\m��,^2�����#D�����_4�"`EJ�I�Z��q'5D���ƃE#���o�1�T��&D�@���L�l����b*�� ��E:��"D��a��l�E��W�B�8�˓D$D�(�Т����ѷ.�$U�N����=D���ԄL�i\Pĸ��
�
�8j�� D������v0�d3&I4Ywt�J�N2D�����U��<ӆ%O>0b�6"?D�L��T<Z]����	Ϳq��=D�d;@�7*~pqH�I�2!Ȉ�U�6D���a��#'��[�ƖKU���v1D�4��O�%A�����!v�vY2� =D��(A *|���B��&K�D1�P.;D��J�K�#>]rl�ݾs���R�:D���`�5h��[qJ���dK+D�(��DS&'��Z������� @+D�Hz"��\�x��E	aL��І(.D��P�&E��[���'Y�r-��/D���v�M�
H#�W9/.JE��*O�]�R!]_7� �J���p�z�"O�� ��E�,>̹s���}�q"O�ʐ��:@�֭ԫ	C�8��V"O�	;��� Ϫ8�e%�)3{�!�"O��ؠj\e|�!o7�4��"OY���4o�xs6͎7<ȩ�T"O���Z�R�H�C��ԣD7��"O��	(�z�QL��p16m�q"O�U��&E$ym�|)�#�r
P�sb"O(�	�ݦw�~1�$�-nq�l�w"O��i'HV�-2�(���~}H�p"O @�p�םl�ְ���E�*���"O�T�	_X�DSaě�
�4��"O�i��Z�F!�E���ȱ�b"O�@&H����0��:B䞼� "Ox���j��^9Ι����T�H̙�"O(��▎n�nE����Fv�� "ONP�w���XA��'
*����"O�r�t�J�٦���}����"O�uك�Vm�@fR�6�$�)�"O� z����k��ѓE��u���&"O�q�5&�,)
�(��_�CV��"Oj4���8Px*!�fH���"O2, �k|��)R�`X#P�T�:�"O2<[
��4�L�z@��i�պW"Ov]02 �+(Y�y����}L�|0"O�xhd*/Fu.I�r�?(D�hS�"Oj�P���G�l� SEA�\ZMk5"O0}0Ǒ)���8���+y)a�"O���ǀG�e5�h�C&!8$@`�"O�eC�a�#W�����.��X
�TBe"Ok1(S���;��ӌ"�Х"O�Dc�E@\�\�aW͔�Ę�C"OnU����+|��qm��m��HG"O����jĚG� aC,�a��K�"O�p��!iXd	ಭ֔`�����"O4D2�l�*P],T{bN��Hݘ��u"One� `X�f�8Q�Cc�V�,(Z�"O�6,�LT,2R�n�29(a"OP�yØ;<�$=�� gp��"O���S(�5S퐶�A�=b.U��"O�1Y��ߣ]mv]z�E�M����"O��Wԑat����+%O܄��"O�y3�GM >�ʀ�`�_��D��"O�=[�G�,�|��G+ 1���[�"O�)�G�W���,I�
����"O�T�Q&A�B���-gdQq2"O��r�HΏg#V�ɕc��UYq"O����n��)d��A"O�zC��	e����LN.r�l��"OD	�f�7" � �*T�q #u"O"ᗆ�@;DDrv�HT8����"O��#��#;�~͡d��UI���"O�� ���q��3D�H�U��L�"O�QڱJ�xG ��Ղ����"O�`F��{�nT8��ވ?�|���"O���@��4x�q�f�@�E����r"O��R� ��>|zIPQ�"$�r%J�"Ot���|Pf�y����sI8D�"O�Z`�3O��1�%�1G�p8"O"܃�+�)d���8DJ!Gmk1"O��B��P�Y��{��M�e#̰�y�b��R�Y;�#P,a'��"ӏ�y�m��~x�I�)�)<��1p#�1�y2�Mw/�탳��]��4I����y��ѼNF��K�Ui"����ٹ�y�c��6}��G�Kר5�W���ybh{�% �~�(���L8�yr�U19dV� ��q��G��y�攋�a�S�V�n!�P���G��y�B	P�b<2S�U`JZ@ʑd���y�I��ocD(K��E��&93����yR̍e��i�&�,`���?�y��Q�V�nqЏ	��VH�kO��yB/�}M�5�t �Y¯4�y�"ض{D^ec���4[IȔA� ��y�O�N&(�R�$Y۸}H�`��y�!F v�k�J�)L��mr؃�yb� +��q��h��J�l�9�Y��ybh�93-��{	 ��2m��y��X����CoRݹ����'�n�sgc��L�����7=z��yI>��ATDzc����.�cs��]�<���٘S��:���fD�dÇE�b�<��)0'�n8s�����)B��W�<� D��&�R�8����0�kxв�"OV����Y�0nJp��bH�`�-!3"O��z����Gz�5B �¤lO>��5"OR(BW�H4<�2��cb�>I^y�"O�5��M �XSs��/ʅ�s"O��	�u~*���/�5p�lHp"OVIXh*�E�E�`� �J|�<��D"<�& ��7��T�l���ȓ�V�ӂțK9���/�	h����VM�え'9Yl�1eW9�M��V͖�)�O�"���2�G�S�&T��#�$�¬G(\j��H�����v�a�.ָB!�`�@��:̄�!�}q���0g^�Hz���*����<������x� ���\�H�,h��,�EA��:��q�A��~nX,���ʷ�^ )E��v��1G�d��ȓ{6&�H���x�� � �Z��̄ȓ&zĸ�3y̌���*âB�@l��7
�<87팾y��­�\ن�k/�aa���**��,؀B�eP�4�ȓO�����ľ;��{ǪA/U"8�ȓtrq"�BC�K��s"�ٷ��,��e60�rCƓ�V�X�4��I��a�ȓ7�l���@��:�l� �.qL���w������+���	��F)Del���[��U��,�L�ad�է>�q�����Vp6d2���d(���K�<1v*�4��{�Np|�����l�<�%�ߠ]*����b8T�^�Y��D�<��h�r0�g�dvt��'v�<�W4�́�	�&�t�@��s�<���/���S&��t�`��pI�o�<��5?<�q�kK�"AQ@�<����8i� ��x5\�# Fy�<�Q�K9A���!� 8.7����x�<10)I�(�T�ÌcQ�4X�fv�<���QP` +�ˎ3,)6��%�Cx�<�� �$j�"\�V��(xd���F/6D�l�S��
��e�+�j�Ld���1D�Dj��
�+��p��l���0�4D�䩀�ֈD�,1*��K.2���v�2D�Z-B]�RT_�C;`Iq��1D�pa�E�G��M�D���-/bh�D*D��;V����:�D�Z����(D�$bq�\�/�r�k��2*$�e<D��aP��uL�H.*Q ��:D���%���
�z`A	�+��!�$����W�]$B�ʤ�	�!�ܢEA����#\��)S#�/8�!�D@��DR���3�.]y���m�!򤏓x�F��X���0#�R�b�!�$�(x*�!��H�@�f�#&g��h�!��,,���D����:C�!��|����I�w�h���W��!�(A^��F��J�$D� '6y!��1>���)�R��A0{!��\�!�>�apX?E�`�H5�y[!���:�2�J���8 ��d�Lͩ	�!�DRG�6���fE�z�p"ل�!�d�0v��	Bˍc]䥘���!�d�U7h�s3�ХyC�\˦�T)L!�d�=K��ƭ�T38m0咱�!��`cf-�/�y!���S��!�� �U�lܳ\Bɓ�	wH��"OФ�䊆m�s�F�W�4�"OD@V�#
|�3�$�1G&�x�"O�D ��ʯF \�EQ�@�%Qr"O�|2�X�P�E��	i�"O�@h ��X%���H:d�� �"O��a �I�?0@� �HU��pP"O��3Ɍ�_�&����!Y��I��"O8�',0�|C"(G�\���"OHب�J�.!q�\�0a�(��� �"O���Vk�/GY�3TIο
�6D��"O�%�`��rs�@�R��OS���C"O4��'O�7�a��GM�@.�;�"O�+��C�n�l`BG^�P�LPF"O8)�F��+:��Ѥ�	)nP�X��"O�h��$;��p���۰P٤L��"On�!�"Z�^P\����(Lo`���"O<� �
�w��m�0 $]g���w"O���� �J���A�@JT@1c"O�� 5byj�	q��R�F"O�S��Ft�WA�i��]�'"O6\�sE�?t�����:߄�)�"O|U`�aR=S��Ro[�-�l-���d;�S���?
��db��+P�Ne�%�R�
�!�d������'@*Z�| �Q�T�!��ËK`���+�}Ԣ��$�$�!�d�	t��0P��= f��=k!�?Z���@) <\v��C�B$Y�!� 0��br��._Z�9S�M�!�dL�Qa&�0(��X��Ay��[%{�!��D�?خ�	�K�' Ϟ[���A�!�dׯI=Zx����0��c`�j�!�d�wAR}��O�x߾�@��!� x��C��@��B|H�O0O�!�$�<�Qc-��<����!�ā�3�!�hs��xt �x!����t�2��3��QSq�هc�!������Q�ߌW�B8����P!��[��e�U�޾�M4��#m!��w� 3�	!BR�JgBE�!��F�\A�0x a΍�,�ء��05�!�D�4"��Q��'�^-!�m�h�!򄇤o�l�g�%pLm��� m�!�$N�?�n=�3/V4�
XF�!�ĩ]Z�H+��m ��s)�JT!�$,�����F�b�;iP�8!�Dؽt����Sˏ=20dS���d&!�d͏E����g��$"�<T92�A�d�!�Ds+F��/�PjHqq���B�!�D�p��ؤ�B$-��3�a¤I�!��B�`�P�Y�Al9)��=�!�>��Yb�Q�&@��ل��r�!�H�TK�Q��✗P2`Lb���;'�!�/s�ӡ�9R�p�N�)�!�DQ��� �`��(�,s�g[�O!��߱"!��jӯ#r�ܝ�f�-Q�!�	4n�jM���5�eJ�]�!򄆉R~�|�Wa,G�DL"0�C2T�!�D[/~�.e�V��i�
x�$�Q'3�!��>P$5ZP%�>�H۠��O!�d	)xLm�Ge���@�%�M,(6!�d�3kRQ�E\Q��yٶ�;�!��L""��tJ������%9��U'+U!���v�M)�Bq<����qP!�� �"��I0>w$���� :��)��"O��c��Ul�e��猜�|E"Oh�h�!��F�T0h�M�q~tL	7"O��R�6*<
\8%C�No�E��"O�IB".�")H�Õ�O�qz�D�s"O-@�GP4|z�H ��{s���7"O��;�KH�oS�XzSOލb2͸$"O�b��?e�����?;���p"O��ZT��P�12w�ԯC�Αr�"O�<�e��(R\����&��"O*|؃"C�*���Y���PY��(�"O��ʡǞ�N��,)tkŚ.��jV"O8Ց��ԶD6���`I�,%�N|Q"ON�J��U�-}��V�&�yu"O�x��'�-'���Y�효U�>I¤"O�婄G�;^��E`�����8C"O�E+���]��0p�aA+U�<)�g"O�e��F\}��o�mw�T��"O(RA-�_v��߭N���"O��%'�.��aϪ\�X�qd"O�yC����ʴ��t�R�"O�	�����*�lh2BJr<#@"O$�`L�g-ֈ:V�`��}��"Ov X�Oӵ@{n� f�J&{8*4�p"Oh=����,���0#)�`Ҵ8� "O��bE�1T*B����	em���$"OĴ��B�6:|�c��c�(Ib"O:���&Y<ZS6�S�(<[���R"O���"�"}�Nu����qSR���"O,\�f�	E��k�=kR��B"O��;#c�	�a3j[�dI$���"O54�� ,"� 3�bHB9�E9"O8�c��@�����	N>nYb�"O�$P��ʋS�J�;Fg8VD�2"O��H�?D�I�{� K"O���	6A!���w�^��.t3S"O�YBe�O�:7��x��@®ɡ�"O��@ulN�Z3bh�s����Y�"ORd
w-M!I�T�G��`�
���"O�aqa��;$�	T D �� ��"OJ��b��=�K��V�4l]��"OR���O�C����"MW�.��""O$�+�HNn�Y���G ."����"O�Q�����Dk��}9)�D"O4e�u�#kV��!���08ht0"O��9�h�K) ��!��7e��"O0�!���!@������M:Y��"O��Y�MʤOS6�J���ъ�b�"O�[����q&<��,2�"O 	&b^�<"@���5~�~q�@"O
<z��T� ��Kf���9�"O3d�H�_�N���/V0�"Opm��CD:P�]d�ń)��"O(E8� ��[�j�F��l���A"O�Aȑ�_�16��0�Ԏ'Ԗ�p"O�E�W�J>��\A�g9v�@��"O�e�Drhb�{e�D�<����"O�����C<�X�R��+_����5"O:%+B�b� @�]�z!k�Ɉx�<I��<XQ�1�r� ��Ě�,�v�<y�'ρ^A*�0�@�w�ƄJ�l�r�<i��
���+�ꌊ=��t�Xi�<�TG�#q\��3`��I�����h�<����K5�`�chC�@�(HH��Gb�<� H-�fH&�����=W&D��"O��V�^kn6x[�B>88D�J�"Ox��r"��iz�$"Bh);^�[ "O���A�խ $��rfX�	��P"OZ�#����D�T��[����"O<r�	U+6Ğ��A'�)e�X�"Oz��tH� r��G��%k�a�$"O��G��=L�~�:�KW���kE"O�j
��m�(��׹m���"A"On���ͅ�),�Lra�2~����B"O��xa�3s�4 �%/��(���8�"O<91��Ϙ���OĲj
��t"O��s,�1(p	H��Cd@P�"O,���i��b��A�X�FK����"O,q���h^I�L�W�"�""O]�B��'?�m[��*r��"O�qs�K�#? ��jZ#]�ݫG"OFiʤO��F� ��*�,i\1��"O:�cg�Y09j4�b�I��R^��1"OR��2�ѯT��Z)9��)Q"O�}Pv͇�u�������|"�)�"O25���^�b|9 ŅM�8ZU�S"O¥�e�ˬNkb���N;��"O\̂�O�/O���#�-\e*��"�"Oʁ�D��M�4H3�LJ#hmط"O�Y���,cN��B  �dk�"O`m��)=�<�7j�� 
�]X�"O �S���9PPf��
v��Mۧ"O�Y��$�#%@ʝ����M���)"O�̉�=p��]�PF\!��K""O�(��IаhT��k�/�4Y��"OP��,T3gx�h֮�sуp"OD�꤭A�f�Z�a荳�.��C"O�x��G]�o��(�vF̸{��p81"O��*Ǧ�`zH:�ņ}�*�˗"O(�X��]�|t����x�p�"O����m�l(8$#Fv��"O��YT�GX���GOžz��ĉ�"ON!RP*:�T���~�ڂ"O0�a6��D܌�"��W!}>�M3t"OH�i�B�d#��vl57B!H"O�����a��q��*S:\.�i�"O��x��U�mpL5��4=��{�"O�IH2EҶ(�
0��뛥sbxB'"O����[����Y;e���%"O|e�� ��t��T�=Ih��R"Ob�2DO�jO���Lv*0�0�"ON(��Z�:˰�Pp�J�XZp)�"O�\�G`P�P1T�@�{l��S"O�]�%eʱ0^,�)rO�at�e�T"O|A��CV2b�HqnzO.Y��"O� +C��O���� ˞'E01r"O.!� E5Sdd�f�S�:P]��"O�����$���س��b��ة�"O�l����lQ��f�:;��80"O!���O�"8���f];H�p�"O��@T�ҙY�[wE#7��YB"O����[f�킥�,>􄈶"O.U��P����B�Ó2T��B�"O.����? ��h�	:,?<z"O�9
%H�1d��li��L��Zt�"OFI�Cg�m(��p�)�;Y�6��f"O>�!�A�$�;��3d�`�3"O��p��zC��##��K�4�s"O� ��20��)*�@�Rv�~�i@"O�@�v�ٍvql(��?\�n���"O����(��y�b,3�`I����B�"OrY����+��a����f=��"Od!ZK@�Hv���X -���"O�u*'�5�4�)w�A>w!��	�"O����Ꞑ�^�:���(���"s"O6 �B���1��XK�%MC2=�f"Oՠ�,�?rr����J�x?,��"O�p��FƱ{Jf=Z��¥�jtZ "Oxu�a㍤2�1���f`1"OB��.�	��̀�+�έ�s"O�m��(����US*�0eR�"Ov����>MK��Q��4E�``�<ApjJ<�	�3��X���uk@�<F+-[pԅ{��ؤ�ִ���y�<QD��9��܊�(m	z|{F��w�<!C�Y�yR8�"b]�v�:����p�<yt%��6]2��5��%r�����Cm�<)0���_	�9[w+� #F1���c�<I"��T�"�$���+`��90�QD�<)3�C�
�Rh;�`�",�!R��d�<�'��H����@�p��ҲF�a�<��(���-1��9�|�Bu�a�<��X�~a��Ö-[�]b"С�$�X�<aǀ�y��آ)��a��!n\}�<�� ��+(Y�ӄ6� �x1@d�<9`�5B��My�#�8D7đ��f�_�<��A�(
n:�5+ǚ�屆�P�<Q����K%�2��q/KM�<q��M>�"���d�M���q��Q�<�r��c3�=b�͏k�I1��ZV�<���ټ6D��$o�Ai��0'�NR�<��Cȴ�N8��k�=�������b�<٣�B߲�
�&�w��QîH�<9a�ǘ2�H���rT2��I�B�<`͖�M�V�A�#��v@a0��[x�<Y&��[tP!j�bPB�ɋ�C�p�<�#�_,g2���pJ�O2h�SMU�<� �sٌQb�!
�>.�!��C�G�<�.A+Tbiѷ�!f�d��s�L]�<YvΛ�]ׂ�a��|��@D�<ŊE�Q�>�T�݀i���(c��K�<1��0j\Y�c�>^��M�'i |�<�s,I0I�����L���ۅn�{�<�t�(g��RH�8Cf�ہ+�v�<!��{-.���R7xa���r�<���@/>��0���D��0"C�<Is�F�B�"E2�O�2j�D�X�S{�<���+H,T[�aY�%�,H�w��y�<Ѷ��5E8���d*��ah��@�<�f�0u|���&�;�2) ��G�<��F��_�8�i�o�*p�p�Ϗ]�<U	W�K&Đ�'_�l�u�OE�<���.���%��+Smi�<��@2$��t�A%��O�T��&|�<a%7JbR,�Ο-��9��@a�<х�4el�sV�5�,!���f�<��j�f"�(4 ��)�h�a�<GJ�zL��0A�^�a�π`�<��(j�.��&,�O�$iA��
G�<ђ��h�¹#�NJ� 3@a�b��<aw��ZVp�!��ĞP�����U�<��O�Rf��iD*�z���UA�e�<� �\�"�(\�$ ��+�8'�!�D"O�T��$S ��Ɖ��LĢ�"O�dqd)�;u��c��a�&$bU"O�@U	[�7K�B��B���CB"O�y���q��i��j�i�x��"O�L��Ы�Jc>����O@@!�D�[�b	n'����B�!���s��9���g,� �!�øZ�p�h�M����(ذ�!��	�r�ҝ��_�NBB��52!�d�dr�`G�-�$ HT2P�!�]�1Lve�t�2_��)�#J�5!�$;BFĬ�%[e�¨�7#O�"����'R�Ի��˨>v9ra)߰�y"�X�c��t�ԤH�p6*݉���>�y"I��x_�i��]#o���@A��y��ʹ<���ߚn&�Q�CH�y�ΨڠQy�X,b.h�9�#�y�'�/���y%�N�R̦$��GW�yBCP>zڰ��v�Y<7�R��g߳�y��ؿhafH��E�65�����N��y�#U9`�t0����[bTR��B�y���1D6HR���8[��a˥`��ybK��O����T>Oe�Y$��y�j�']oҬ����K�f�C:�y��\JxB�nS�z�����yR�5[�~�0t�X�H�p�iG���y�jG�`��(���q�nM���M��y2��z����1l�$_W��9��U��yBG�; 	�M�e�I�D�T�2%��y�-�_�XytEX�B@V<uIñ�y"&����$�*;��,�A�	"�y��@0rK�� �	�<7�M�B��y�aL1A9�l�B�$5DI�`cA��y"�M�'����'�(ľl���C��y�c�8�(A�	�$ �ۣ�)�y�G΢�n� ËU�'�KS��.�y2��9��ڎ3$�`�5�*4����'���tI��M�)��$�.���+�'�b������$��6�l�'��A�>f��	;��${;�HY�'��EЗ���S�BL���?w�
]�	�'J&����nG�ɑr��g��+�'�6}���ŝPT�ar�[5
�����'un8rM�4����)��z�	�'}ʘ7��� �h�\<�RĠ�'D�D����,x��$�^8}W y��',�|鐃��T���de��sc��(�'��6��.�´Z�"ۧg}�\h�'FJ�C�\+`C	h�I[3X��x
�'{N0*C�N�����!aӥI:.T�	�'�p%	Ba��yq
B�4<�k�'��-��O�S�a������'�6 ��iX5&��`�oT>i�d*�'�	�"*�
c����a�D��'tၤG��Sa@ċWT(��h��'?�}ˆ+ƎO7^Hr����'g�h�
�'��ڥE�!J�n�fG����'��� ŏ�K�������`��QA	�'�1� J��K�H-6���Xj�!R�'� ��爏7q"d�j8��'T���RD��r��9��L8�l]�
�'�(�1�g�>.O8�Ԍ	���j�'v�d.[/`�N��L��yP������ ���)s��q�Bk x�j�*�"O<��L�8��u��0�T-Ip"O�H��g[�R��A��������a�<�G�J��$�ק�7__<���V�<��B�j0h�E�L0B>�=��ACS�'+� r;�@lZ\�'38~�1��Ѥ>���J��F:���=�����2��f�p��'�����k>�)�ix���VԻrq0�Q'�#�u�ە%�$;���*�l�8�j G�:zfi��J�p������%.#�ળA�MϱO�d���'����i�z�B�6f0Ҥ)G3�����OP�O����O�tP� ݎ|�$��G)W�M�: �'��6��O>6��$J���a�Ş�Vx �b�)H�Jn��@U�v�n��x����7��@�Z�B��B"�q:t9��P�4Y`��+ )J�*T�	�V��9�c<m�q� ��w��WcO#D��[w��)~�8H�ܴ`��xh��W�F�P�2�)�9�1:ԨFq�lA ���\c�`Lk�,����
�@AX��4h�=����H (O��џ8��f-��ԭA�G�ZPV}d���d���O|�OR"?�!�_$uP��(Z�f��!!��'46��O��Dئ�O3��(=x�lӕFݏb����{���D��З�i!ay���X馍�RCϫ(鶑���	�T���i�'+W(���� [T����⟤�É���D^��*�[�Cn����o�3�U�w�۲>x�k�۪]���"#V?Y��k�8'��]��OX�9�%΍N�`)�.:�aƎݟ���$�Ɵ �	`���<i����VIk���%��:q:�=����O�Q�@��	gu�$���.(I����e�?NK���!�i��6M*����>��<9q��f}�L�a� � '��	��V���?	���?�u.L����?��	J�m�Ġ̄K}��F/��MF� B�Kܭ;�ɓ�]����
� �#?���R Pb<h����,{����F_�H��!�sլ�k1��#l<�և�|�]��Ͽ�?�ߴ-e������+L���q)
�]�9�r�|2�'[�T>1#`�?;&�R��%���	t�9�I�=�#<%?�{3L�;d����Δ�L��$j�4�?�(O�9QDQ��M��H���z���OY3+��+�ME#����"8�*|9�! M�>͈���YH�c�:��hx"2s�zy��@	�Ʊ�q鉜j7�T"!�'E�b�y�-H�v�U��B��'���3��Ѧh��ܻ��6��Uk�-�`��k��e�IƟ��ߴ�?��.��Ђ��[nT@p� �uc�ҁ�	/H��'��iݽD��A}�B�7��4�e�_
V�8D��	�9��ߦ����D�������8�6��C�Λ����[�*��?���G�ژ�?���MC��-M6�R��0@�rT(��V-4��<���9$�"wK&�����MB�+���	s�)х�ӑR���蘩neZ�ĭ���CqMb]Zٚ�+� ��q21�[�#��T(�=���>�!!��gJ�Dx��N�/�,\�i%��9���?��iU�s�Z�b���S�0���b[5E�ƈ��O��d.|OR7����*a�Ӑe
�`�F�\Q�Ԫ�4�?�M>����M�0%�8i�)�`�T?��l��j[
!��՟L��	�p   �   ,   �L#�靱I�ƹ�tC�&�L�:�.ħ�~��w�P��A�N�Q��P�F�XECDߦ5J۴q�`��� �,_�\�ퟌ9�@��Ŀi�06��֦����x3��3IT��3�c�j��8B�KH�'�މFx�Ħ�JE��R54�B��Fh�Hh��<A�N>"/�)�ae~�i]�mD��m������-Xu���o�LZ���`X��烈��M{��'����ɛ���#�y��	�3F�A&̀/�|d�aDZ>�"� �d=�ap቟ ��ϫrP\�ˌ"&Xl�b��S�|��'�l\Ex2�Tr�I�3��9��~RR@Q�k�=@z扯#�� ���	
 s�!���v��cCI�DG������O���O�l��$��;/^�&�˽+�l��Ӝ>��+�(>B����dZ�+��˷n�e6�T��"{�hM���-�O
Y�b�Z@��1��j�J��gӱO���Ĉ<��D¸e�X�`ǋ	�nٱ�i� (��I"/���K�d�l��T(@Mڜk�~�P��F�1��d��O�����F5�U-֖5$
��]�=�<�L)�;�hO�QhY�}�ָI��u^DA6�O�s����!��'�DI!$�����=Mhr(�'�"��Nqy���_�F�+��������Cퟴ�L�7CQ��랅Z���f9���Sr�>I�*� ���i�`	<�$�����x}2K�T�'ifUFx�BM��Kf�Z�ag�(�����y�K�$8 d  ��: �>@�����6Hj�g�aM$x�G��O��$�O6�DF�����?	�O]Z��ڴ{� A�0Ώ>��	樈���L��I
^��7�R�d�����"tR~�9fnZ.`�ar�ץ�MK'd\9���'�׌v��`$
�tH!�E3
̽0ԏ�Z'^������!�$�y���DDڍm�δ�����sR�d$�OJY��JYɦ��	���mک}/�Q���	W�,�2w"Ϩ�l�Z�$a����?���}l^�H��i�1O�n�;p%h)�r�@2|vD��!�����J�m�O�O�!`Ub)(?l)hv��QJX��d�����'M�O]ȹ+&�~�!J�烧��L����O��:�)ڧ�0�*B.<���Af3�ܐ��I��~"e�:P6h���
OD�ʲ@�4R��L<��i���'J哠O� �I���� �S?/F�*���,>������?q�����?�y*��'Ő5���8>�H�sB�w����ONM��)ҧj����Z�Xa&9�V��,l��'�2�*�����H�|�qD�m%P0p��*g�6�:�"O��U��v�z$��$W�R�h!q�I�����qr��Oyʜѐ�Ӧ:�P��g��؟��	͟��#�r�����	ڟ��_wd�����g��Ԃ�,]2k@6��"�Ϥ��E�^�1ד3���5�̹�}Ek�,3;�'����b��,8@f*Y
�R9� �ނ��D�*:�����O&���O�7�� /�J��N7;��P� ��!�$�>,D�Lv�4�
PnC-���I�����<ɡ�����uREE�~�8u�C#U�L".�P*A��?����?I����O���e>��ӎk��u��	=��Rf�Z���3��'��q�ݴO�,4I�C/��I�*I�Z���*?��7m�>v���{���M4Qx�#�Ȃ��xB��'�^uJ�A�'ޭ(u��yb�S,pVn���"�t��D����ɉ��'��ZU��>���M{��L�wy���r�KTF��2O��7lf�#,&B�'��ǆ�M�ÃDG91�(��m ���wc]�)&ⱳÎ�U��;��}�'�\�x�I��A�0����	b4M�S���Cw�K�4QT��N��~5�#?�G�O��$(�	��1�1A�ΰ �\���U���>� ��A$�.��\)����n	�'}����
a�a�
��2|2��]�|n�x(*Oz���OΦ��	՟T�O�@�5�'�v�C0P����?�0�sٌ���<���-�|&� �$䉲R
&�x�+0U갘���>i�O�b��H���bI�/$xhH��^߲�X \�`���O�b�"}z���)7�A�sDF7��8됉_l�<� o��[����p���x��@h`	k�'��~�ҍF�R�P$0q圄%T`�%O$+���'b����*���'�r�'2�qo�1&" �Y�J��6��h�)8a���'l)�S�\2Q�X���
���X�k�g�4�{�g�2�M��V��yTM�<lJt�,��Đ�0a��ѧ̷9�t�h !նa��4�?���?��S�Y���	�����L$DB��"N��� �7m��0��ɍR���lЇv5��yc$K�TꓙM�C�im1O�SyyRDѦ6�,H*�����X���\�V�����rm��'���'�.ٟ֝D���|b�mF릹H�IBA�`��+VR|���4�O���M�"DK�" � e�g<��"���I؟��h�L�A��H�[F�@��mÕk4&�(���ZH<Y�#R�:�`��Ŏ�W�\���C�<���� �\��쟺hEtLY2���$@�o��Y��iC��'<�F�	�+�䱻0�I3kB���ҩHa���D�=w���D�OJ����>�$(�i��k%'Y�7�ތHE��A�6���b+���(D��J�1
��
� �?� �C$͒���O�Y8`�'K�����~8.�#%�E%?Ep�£��v�n�$�OF⟢}J"��M��C#��ﲐc(�y���q�'��E�E匢6 ��
$i��ɠgo�<i#���*��f�'�R>�9�b����o�/��ؐ`��fA��g�������1FhhK�����|r�\(<ۂ�@�ZTz�H���+��zc�"}�-Xp�^(�u���|BS��@}��ɮ�?��y��	Ʈ,fƌ�,X�R�\������!�$_	D���@"˧02��Z�ė_�Q�h���)�7�
� 䟈 �JT:�E��L��-�������6BR �z�$����П(�	 �u�i�ll��V$En�=GLۀrĺ��M<A��o؞p�����B�d̫&��i`�ܙ�f1� n�a{�$�;)���rLB�4�\s��[���m�T��tX���V���"�>tx� 
$r��@.D���s͘�����6�H
w��Ĺ����SDoz�4G�-�F�"uc��po&��'+�U����I��������\w2��'�IV�J"��n<0*����Ȧ$κ)�Ǥ�ٰ?	���9���L4xm��ڔM� 8��-��A'�O0�pd�i�r|�f�C�uTIc�J�s �r(&$� s��Y>��<]c�IHv#6D���f���_]�a� ` �?���0 }��?�ɚ���ߴ�?���M#��/V�lr0�̼~��(���D92�bD���'���ʷ9#�|��@`vȢ������\�>},F~bgڥ�LY���F��%���r�c!%�(�n0���Q+3��0�T�I�)2���O�mZß���)��@��]��l����8q�	���?���'�$�넬Їc}��£/��Pi8��ċަao�/:�`Y�RdQ2��������.r��/O�cE�æY��ӟH�O�pt0u�'|�� %(+� j�FA��XIf��y �$�1Q��d/�|&���w��:|�5���19њE����>�Q*u��H���Q�G�� �� `�7�v��]��V��Ob�"}b��̊�L��,�:�*��AEX�<aD�P@>)�3cW!So�ٵ��'[��~�G�\���8�G��?��!�D��~���'>b
e�����'���'�b�s�Un�
z3�U��!R�y܊490mȹ.��O<�p�旉��<I��0P͈Б�A�x����%��H�	:��	���'W(eۡ,^�Zϛ	�Ĝ2sE1?����)����?���M��f2_R�	Eb�=w���W�<�����^h�$�欟�Ky����d�R?���)�I<��#.���,B�}�.9�`FM�<�r�&c\蕂�<:�L᠀c(<���5&�ʵ(�O�n�u���	�W0�B��*,��J䅐!W׆=��hD�cr�B�	(_~��[���h�zA�å[(BB�)� ֘�&�K�/��z2
�;��"OԼ""̌3Ȭ�RS��V�lI�"O��p`�5�ZD�%e�5y�`;�"O�[7�ı	�4q�!�׾���`�"O������P]!�l�=�ʨR`"O%�F �}4i1"l�(��ȓ1
r@��ŗ��b����>��I�ȓ2�^m1,B����A֭	�@9��fƄy��3I"G�^!X<�ȓg
Qx@�6E�yr
]�XgD\��j����J�
epHq�ſ'
Մ�U�}���L,zQ&餦 f�|��,��V��@�P�皋x�&��s�E�Pt����o�X��хȓ;~���P6m��Չ��D.b�`�ȓ蔘��ʋ�{���N�=a�%��n8~���  *R��XЎX�T��\�ȓt�� G@6C*��b֘.�� ��my�W��}��Y�EnO�\)���ȓ�Ń�ϋ:	|a�5�}vޜ��fw(M!d� (�b1����:V��$��W��Q2�䁛Z���w��4:���ȓ4�T��K��=�8e���q�����A| ����%K�4u��iƅ;5�%�ȓ.^�� � 8�F�������d���o��g@�z�NЊ���{�2�ȓ���%.��|9��*��C=I��GЌ�y@ND/4!��-�6!���>
������";}�t�A�E
[�*��ȓqXhEy�戊*$� �'�-�>l��d�Pd'��R6�X��O q;����T$طb��z�!�.V����6	�x �i+Ŏ�C���C�PY�ȓH��$�jO�.|sTf�j�����U^	s�E�7'bP3.8'M@a��VP��a���O�����%�7f�\���[YrpN� 5���@�D;]�5��|��}H�eށ'���C����A�ȓ\��ұ%�6*�(X��ӮDB,���0�V�9Vj �l���rE�c�\t�ȓh� ŋ�s�I�!�ީa����ȓE��=KO��%Zu&R�d��ȓ&�S��H=n\�1+�"j�чȓB. u�q$�����4Dd D��	?��ASTV��Z��A�����&M	�ʀ0Q�>D��j��ٛh��p*`��t� �V�1�I ��J$�MV�O����V�M!<NR�br��
�� ��'YNP:A`)�9c���<��3��$���J��7�<q��H�"���f�;l�3 Y�<��B}���a�?W�EC��óa�tat�Q	\>���IuڀY-U$s���`��%�$���\�n'�QB��	5�y"�˧S�|�!°d�a���%�y��ˁB�U�R�B*�:�H��"��'�`8�C���kX4D�&��#v���E�z6�'���y"탺f�"zs�̫8���B �Z�&��ɒ���	�T�Q>˓�(���OF�o�.	�weC�bi���V���Ӳ�ܹ1�R�Ke�62�cE��=)�ص[�y�X���+W���E�"d˼��5\Oh`9���l�
5K�'��\��g�N\!P�k�/^���'��A91m�>
,]�P�L*M��}��}�
Ӵ���.*�'s�I3E�ڋ_8�}� �'a"BĆȓQj�1ÕO�V�^������}�ʬ
���3]�qOT�}�Dn8��B��,_zI�	@w����@`���k7E��Ę+.�@��S�? t��ҡG�0�p���:Q%��"OFH5K�`�Ъ���F���0v"O`�yB��w�ԣ2j���l�ֶiN\� N\�S��M3�+�>��)��#؃�<��WN�W�<')�-3�FE�e$(Fd銣��M?���*�(I9
ۓ[Ŧyñ�PXd�!�E�*�x��I�-�Xe�����cҼe��K�Mn.��n�x�@�k'D��{�����,�zl�1N��g�"<a�!�т��7r��|RN,lh��%�O�H����WS�<�w惠Z��0@�`�+!�rxB���{b0 �5Ό��ҧ���C�S%�с���`���$Vl�!�$�2A�-b�,ٓ_\��慛�x��$��UǊ�Q%ř�p=9�'Иk���(�'�z_�A��Y��ӲN�-.�� �3(�>n���b���-���sV���r�����j���s�_��r
�^�*�;O*�t��N8b��=0@���#�ع�M|2���^IĔ{�A,��� ��]�<�!��=��k\+.�򸲢@�n�*D �\h�̭����)iE��'/@����:[T8��uˑ3O�dI��'�bÜ3��DoK66͊�n����c�Ò�[��}�FbC�\Y��	K�J�v*ޞF�� `m��L�@���Z,���"1��z]Xݒ�b���Eu�2M����J�z("���G_��M�a�(>K4�y"ϝ&S�ax��v�Z�	��LS�d>�Pm�g	P?6'�X;�� $!��ܯ[�L��A��q�T9��W�i ����ԯ���(�Δ�,;va��s������Ҙ��;X,q"+3D����iݙ:��y����'Q��Ԥ,o�ԕ��ކ�p�p�-OG���ɕcQ �(�Iσo3v�c�,? ���DFtJ���g �2+Ũ0�+ܦ�Y�qi\�x�qs�圬0��uґ)1�OV��Z�1��I�a�3-����D
 N��
�H�kx�x�v��z͉O�-�A�ݮd�м;W�ȱu�$�a�'�F(Pv Л�~x�m�/aZ%�(�c�qp��ޢ���2�H��I?��c�ԓB%"ǬC��B�I%=�xJ�kCFa��xPD$��6�ǔL�hQ�a�̟��=i��+6�+��^�������@؞�#���|l@:��'���(�&Hj8D�$��2w�uR�'��(�D�z�(w+��I�5��k�~�~���J /PF�,T���\�!�1����i��a��Ң��+�"OX��AhsE�Y���'��l�T���n�D���Q�J&O��E��O��3���6}����'���"On1��愮$(U���"F�5�P�V�;mJ�B"R$@zZ8RD`�"	@����\i���A �Mj4���i��QNa|���N�@�bPeDL�fƃg�y���NUi�q�Ŷob8��$�q�a�u@�%��<��iR�g4џ4��A�>��Ґ��@��V �#��$q\X���nA��y�-R	2�qb�M�2j��B�ش������2�����)ʧ~����`�����gV9
f6@��j��J���4@��sЭ��_ꌋ6�>��@�%��!O~�=q��+9R���="Ά�1t)�v�'p�=Yr��HyR�Y09�*�����S��}p��E��U�dD\�E�h*�4����ݪ�������M<�X�W&��Q�إ�1�	=|��ќ'dl3�ݫ���wiQ�N9�\��y�c��0� ݪ�GƄa�@�3C���yb��� ��#0���PV��S�` �	"=
�H��Mӳ���g��at�2��ė<Sʡ!��\��&�	�+>�z2/��f��]@�Dʎ]*�@��G�p �u8���R����C��)z�;��م6C��0Ή�?�܆�I�:4�����L��JP��:o`➌˰��6	6�ə�W?b9�b:��Q�Pc���Y�AƮgIp:��Jf���r"O$�8��U��`+�I�@�������0�u�7@�|�Z�Y<� ��0�	ڪ_��׹RPM�2g��<ʠ�F�е�!��	�U�ĩM��z�N+���� .O�ʼ���С���w�]��I�T�,���,p)@���<��$�$"S_����>���b��T��y���8K�@8�%��&�|X�ź�l�Q�\�t$��� ^^:����L�k����C�0ђ�5�w�ɑ1Ԝ0��C�549�A��-[�8�h)s�I \5�x+�'18%�0������s���[���ȓ߼}�6�L�4��a�5�l�ԁ� M�mM�t�I߇^� �&�;۸y$?�f����� ^\r�H��4�Ӄ�؂�LȐ�O��)
W!A ��UK�90�{�+�q�`�`�]˨������gJV'MQ�\#1�U Fʔ��q%ݩb����3�+<O���%\�g��Л�)
7�PI0�N���)��;���3��Q��C�I;gɄq����,9�Y��/\��G�l�q��~�8�z�(��bɘ�;��N�1����k��@�>�r��Ht����"O<�J�G��Mc �s
S/!t���P)�(Pw"���&��u�0�*����s�Hu�u.?���;S802F@&���C�Kf���1��S�nx���#��aO-N��TS�/�1A�ʉ���_�i���d�O�T��x�˄(Z�A* k�0����'ɔĈO|� ��3Mh=;SF�9T�4�2h�T�U
dG�&��2dDO7K�Z�1��%�y�
Q,BD�p�퉔3����¨`Ol��c	�[
�(3�>�j6���;�XA��e@0���2S+(��tIuӼ �R斑b�P���o>F�XF�l��Z~�<Q���1,�B�Q�K�/���1�C��	�Ҏ��F�\]���Ȟ;d�a�0/�F�A�)���ݼ3����m�Yxģ��Z��ђsC]����Ꮢ
H��2-��X����GK� &ʀtB���(����K��|�.P�L�<�
Y����7�"�w�2����z�eS��HM.l#>��Qp���9l(��!�/�u�3��1�0	@6R:ien�á��y��Sa8��&F�`����e�*�,��Ed��t��r�o�Ĺ���_CJ��W�'���U��/�&�Χ~q��h�(�=]\b�@��a����	-�4�A�Vl!�$ 5(�E5�� ��v��F��$�|���ܟ~jH+���l:>xZah
h��͓��\c�,���8�4�! �+s��{��}�4Q8H�WLi���5m�ȼ��N�ֹ��40^l�vMJ���?��q�����'���Xqn�<
h����̃�h$���x�
h�GO�:/�]�7�[	%(b,8GaR)�$��$gx��@��p*����'�X�`"��y���K<B�\PӋ���w�pq�X��~�P����s�k #RL�>Y�Uz�/�[u��+"O|��S#����+��R�=z���p�'4F�9����	���q�SZ�Ф�)Ȣ{��q�؂��Y�ȓL���j��؞F1�	�T����'�0B*Sf���{ש]�%Ҋ@x����6�5�*,D����¥+}����+��Q �(D�X�1�O�sXȁ7�[^@M�@�&D�`�,�+�iZ���� ��d$D�ASĄ�P�Ht�Ҋ#�v8�-.D�$�CS�V�iE⏯kJ�J�*D���G����ë/7D|:�k
��y���}�9�A�O�@�@�<Q���[�fAs�*4�BdD�<����Q��`�g�D�u%$�x�<�G%�`LuC7�H� D�8�,Dy�<I6��%��'�6W}~% rL�<��6,m*9p�E��|hR�\M�<�"�]��z@(��
�]�$<�2�VD�<Ab�F�
ZT�6��h\F�T�D@�<���ґkO�eY��.��ccT~�<� �9lx����L�c	�H���T\�<YqCU�x����O� �	�PZ�<�FL�W��j�8�n�-��<��Π���[�8,A��QW� ]��|hm! nU�M�h,����M-R܅ȓn��XRI�9|i����Q#q�ҵ�ȓ�) �a ;T@�08@�Y�[�؇�,�U����vC�#7��W"��ȓm@�U��䘎'���s7��H�Ф��U�Z䪥j�s��L{f�14%�4��H0*�a�m2:�ȑ�2��+=�����32��A���X\YO��W���9�dd�'

A��l1�b�9b҆��ȓ^ ���%�E�Z�W��P����Q��%�1z^D� �uꨆȓd��̋#nn�`ej�5ĬT��4��Hjb��<�Ղ�!U�*J�ȓ;��IH�"�V?r���K�~�>��S�? f$X#�ʹ7���чo[�9o�d�'
O�iC&D�~w��y�)s��]�Bo��y
R�;�v�� ҟj���Bl���y­͔HL�L���	V8`���镶�y�@�&��i7��H�d�ZD���y�=-܂�@���8@���;��Y�y2��W$"q`��h�@���-�y�l�>��\�c��8
X�y� -��yr
���n�CD@��-kԨ�@nJ0�yF�BF���'	ظ*� =z ��'�yg@0"�u�b�7u�����'�y�C!h{z�3U�*o��H�����yBD�=<� Ո�N�r�
�k�E��y�a4e�rQ#��Y���	�j] �y��,�ʦf�R���Aף[�y��e��!H��>G�j��IM��y�9j�+�+�11b�j�/�0�y��{�� �t�N.!Y&���eI�yR/D��=�B%U���l�� �9�y��(�~u�*ܹ{�0H9��;�y�#��?��꤈Q
#�j9������y�Y,䢼c<x�ā��y��'�Xm��#,�6���� �yB�4��X�n����[ �y���j����n�X�S�D!�y��1� �XPaS�`�\5��E��y�i�� �h XgO
�[�����K�-�yR�R�]N�Jw�R��Ӵe���ybdF�}}�� �����
� > $���'��!��*`q|��J؉(�D�z�'*��qƄٯYi�ݫ�Ȱ����'!�p����6<�k϶E���'h�r�O�9���A��l��}��'��1��DJ,2b���d:w�m��'r��˧��`E����� �h-)�' .s��B,5���4��-�<�j�'.X�A��+��K��N�t$ư[	�'(V�#%iQSOF邓H
*_Z`#�'J��Uʕ�,�&؛���~_"	c�'ؐ���ݥf�قG��*p���'Kn��  9l��rgf͙P�r
�'�n0����5-�� 賃P�Ef�Ȓ	�'8��!�#��B<�9pC&^�7��h1	�'�2��4��#��9#�٪2�	�'��[��h0r	�Qυ<~?�p��'��-���H�P3�._�xN���'�6|h䃋u�F����V}�
�'uj0�E���P�+h �y
�'��k�n	�4H�tqȀDu�'[p�85C,\#���M�{}Z���'��1B�J��m��u+e�@�g�B�'��:�둜?�B�2��>]p>�3�'�:��C�.)���$�G�I��YY�'���RÈP�&������xdI�'�e*��J��0>y"�Хʴh�6Rܮ�q�eIj����M��+CB�I=*HZ�j�)�x��q���O--��C�I�t�٦�g�ʹ��h��p(�"<���r3��y����Z��S��5�j�3 �S�I!��)	�(Ƃ�5XH�9��iZ�BLȽ� N��e$�O?�"Ed	p%�t����N���B�Ij��Ks��"\�������l扸0�
��I�S��X(C�S�̠`Ɖ�?ǖ���%�O��y6D�(%<��� B�v @�"����mSr�:_+!�1kyZAXa�^�?�ʰ�T�͝&l���S�g��F�� j)�*v`�WIX*4�,Ag"OxT���L�/��%��g	*}���Qt�F� �d��{��9Ol�8�ƈ�W/*̲2e��.����q"O��FFL����D
(2����B9O�Ļ7�p>��.[�+���ǜB[Z�l�X�0�R"A�d���S,���U%N���uny!�d�&6��3K�,Kڝ{3��{r��E������ G-�P��d��5�y�%0X���FŢg���h��V�ybD.>��IёCW�Y֌��m��yR�շ���sn�8A�1ȴ���yR옭':
��GH��Vu2�/�yj�rZ������،#U���y�jO�_�b�s@��?nR��!UJD�y�đ0#@���X2i��\����y2LB�KDG)_'(=B�ȓ3_45�t��o9�A%�=�0��Ґ���®dm�d{˟�~J���'"O��q��4y��B��'g���C��'rR *���O�C)�gL{vD`���pf!�K�`�P���yeT=#���G�^sʩxBl/���򙟀�@�V({n�P�$W�Qv��1�J<4�ؘ � l���{3��hǸ����G�IbH7��8xgv�������Wr�|�P�ӳ���&E�1�`�6O~�W���	Z���ƟX��� v֒�I��PJTscjՄqz�`cOl��v�G�N_�e�b'�xp�>��/��$���sY�����[ٟb>M0��  )�8���O9������3D�$B�O��c]r<c�e��0����s�APw�yy�-�f�fH�	�~w�>�Kᖟ�T$��.�򝨐�F<X�`��n2�t(����-��� AfD	H��!釥P�Q����.T�V�����>�
���'h8����'�^အ�7:���*�j���9��J_�q ƣ\%Z�>t�c)�R�P�1Π��V�|B�I� �6� ��Ѐ��ӄd�\�'����#>`H�h�ɆW ��Ş,��d���RA��a���ȓe�@�{�-��2r�aȵg8���'Xrh�$+׹�?����O�'���Jv�Q"a�4jJ�AbFO���	ey��"-O�-��Y�?>$���@�+"l5F���vϖ$|�I0fMPBM�Qa��'�X�S		sl�5���^-l�sL<iF�����	��Op�2î-�P1+����`N�4�c&T
V0T���{U!���U�Be�7�ʌ&iv]�V�.Y�v9YA%D�=��nǵ��'�f5�I�rWp�p��y�}�pfޘEf��c�E�cP��6�8�d:7gF<�4,�#KI�(GBmC��ыl��'ю��I�WY6�*�o���d(��-H�r��+E�P�30�`@� �d}��	���Ћ �����i~Ā`��ߑJ�T���ٳ19�q1J(vj�� �X5=n�<�k�9W#�x"��a�2���	��졶A�)��	p�f��Ge���@�3�'��O�N߲6j�Rp�ޕG��F�C�E(#\c<�0+�,T�]����8=��;�V!H3ҭ�F��ş�яyB�ۧ=!ʩ��% �c~h̻|K�(k�@��B-K!�@����eܔ��[�3o���K	�"őeH!�d�03�d�'À"~4"x�q��1cv(�S���$�5\!&�$�L�,Xh ��L7j��xb샘rA�a��C�r]���I(�Ԩ��f9PI�E�b%�"c��RuF�:N�V���Lm�B	r���*��O��"�����$�����Ř>��Yb� s1�	�A�T��MR�	�`�`A z鋥��2����$�1r2Ȑ`�-�J���;�QR)\�I��
5t��5��#��"���O�Q�'�<�G"��;��}�&ÛF~�!�;0Nf��cd�0$�����ۙ�jy��7���g3l���*��7>h��l�2��A�l�O�x�&; F`��C�8TNF���"��WѾi��`埤��'y،�b�s�!C�,r�e�b.Pk�`Q��K�O<PAC�+8$^ ��D��?�f�8�����dB��<Y�ю<CN���"	k�&%[ǃ���sd��f�
4C��ߠNFD��Q�ڍZ�*�!6\�t0&����	�M���g`��*c�V� ��1Yր�-I.�E �n�bo�����t�#�O��go"����A�Gj�2d�>Pbd�'���	�
��X�g	5���֮c��T\c��b�	�/�&�l lр�H�!*lO�@ -�>a�"'`Y�����*��z�Eʊ,�!Rr�.\�ɨ &�O��:Ċ
e��X�ƭ����'�P�T�^7����k�ZLJM9�}2��V[B)B�:�ܑ!#���0*3�P�G�"� �2� Njlk���!b����#�	S��%���ѐ:���O�Ĕ�[�&߿Y��p8���O)�TX�42���3�L+nv�A�%�n�("�d�OJ���lN+0�B�n(Vг�dGy�������vcNB䉟)��D�Q�+9�\����EN����"V�yEH��1��O<�[f聝-��d�'y\����%��]�p,�ݙ$�2G�B��4Nבz�8�����°2!)\�_,[���m<�ɺ��3�B�yw�؀q����ς�K�.i3'%D�s��-X��D-{�Ș1��+ ��e	qӱOxX��K�40��'k� z�,�d��l�DL�Cۮ4��rp�[}��R�� ��Kg�A	GG���U����=��Mg��(��НcP�T���Zd@�uN��R)�: IU%��੣A4z�t��ɽ#��tQF��޿���+I�\� �^#E8l�P��i�<��cƵ0@F񓒭�y�6l�i�
Jz�\
`/	��M�^�F���k�բ3���,&�Y�i����Ƒj��bM�Bw���)�`~az��[�{�
p���G��U��Aԍ(����&�*N��mb���tY�݋�Ę
]�"����F}��C�M,�Te��@B�4A�$�:���}j��%��8���=꺝CQ��1J��I�FZ���ڡ��)4���*G6(���Yo��Dg� R�l .re���/�O*QSt�G�ou�Ժ�A�g̚\���x��R/X�[�D8s���q�PPr�_���đf�.i��w1V�P�k7p���ͅ�i|���'>�r��ƴ`b��!+_��F���H8G��L�"���$�C!�<�5��X4z���薑Q���v��|P���N��g�_�~v���U���ꓬ�=a��T�g�0o¼��'�.I��x�����?��n����Q�w�.Xd�<��+:�	��)XV-_�y��0Z��\�{  �,�V��@ ���`Eђ*yB�QЏ�M%Z� �����I�NQ=b�x��r�RФ5[aᛸ$m�!҇,*��h��'P�9�N��P��Ňb���m��SL�%btQ.u�^}*�i -�u��"Ѱ�s��c`��� ���S��-d�!�dά�0zVj�5YR4����q"��Dy"jϮ[J 0xRb��R5���31�k에9��ɤ#�0S��q���K)���	'/)��*��y�����N�dH�ա����l��!�S�.;*5:���#���{ +
08�Ȓ0�S�W��OF�Y GG�2�u!���33����d#9�,�ȷ��X�$�F$�9b�f���ӈ�M��b�2d�
�!�(c�AP�!S>�v-Ar�?T���r�A"���#N��%x���9��Cс�IRZ�� J�����AQT�<� ���$�'�*18�I[�C����b@1(���Y�B>D���.
&����\F\X�'�|a�B��N�\p˱iŇ!qRQ�'����k¨K���'�<7�������� ���t�F���L��r�bv�'��-�G�ɭQ� �" G�6L�.)q����I��*��	�A�!��8���)PTpA�-�\P�,����O)�p�B_Ķ��ee�&"�c&��2H�,�Ad[��m�#�J&����2eP� 
�:�A��mh訢�|Q8$�@F���`F턴<�x��y��ڰ~ǄPCE�փ����eW��9"�

J5����I���O��^b�BG B�7� i �H�V�E	3.^>��8C
Ot�G� �	p:�D�R� >RE*H7�X�r�|��P ����'[���A�Z���I�2������'�&ق� !6�&�y�P�<~��3�'E��[��2E ��,	�g%vի�'e�片�FN�ʶ��%3^�	�'�̙.�(��	�*][��'O�@%��3$���
�#�B��'��=S�S�y�&1�R�[�wlX(��'�vM@s��D@�p�Ħw��ɒ�'Q�T	���2�`uA�o4(�{�' & b��ǫeվ�s❪d�<���'�N|�v
B�2R^�i*��` �`�	�'"\�a��
�3�������+��c	�'(��cS.���÷� �r����'8.��ug:Sa�}	���d�fd��'Ψ�c��.'tY�F(�^	�':�{iW-d��U1r�,�֍��'SP����5�y��*�|^Q�'�ޭC��ضkݒ�re��i^�z
�'5�!�#ƝcBhHu��]�4�)�'�nҴ�&�l��o͈R���'P=i��
rՠQ�T�P?P���	�'���J��HC.��A�� J�ش�	�'� ��F�ó
2t)%��3Oƚy��'�֭xN��Z�g	�.�$ ��'�Zi����8y���]�;�x)���� ��òI�?
��DQM�:H4U�E"Oj����[��m0"���I�;D����LvҐ!Sb�9a�	���$D�X1	1%4h��@{�,�%�!D�|R0�{�œ��*xb�C��>D���3ņ�+vt4 2��>I.�&&*D��j7�Y�jb`�&/�58T�7�(D�!��E5|V
�K7��G|��$D��P�,ڮSD�I����0��-�ҭ6D��y�g
�Jp�QD]�P���I6D����G�a�伩T�Dc�Tc!�&D�t�%.�-UGm@�.�vt�#$/D�X�GHC�U{�p����>K�(�	9D�܃�.H:¥W-ȉ,&�kF�8D��P�A�.7b�A�m�6i���ՠ4D���sb�-T�w�9�Lߣ68�X��'�*�+��?q�.��"*�2'�8��'+`��"�*v���z�i�	!Pv\��'�@)�n�M�,P�2���\��'ܾ�q�NM�4wKN�;T��/�h�<	�f��Pע��%A� ��&E�g�<��
F�2۰)����8D8��3 $H�<�b�7Ϧ8r��8���E^A�<����9�b�厏�E8�K���~�<i2��i����Q5~^�	���{�<�p憬O�"qC�-��͂&��y�<Qg��`���� ��"���i�<��E
�D-t���� Nt@|�<Q��@%`Qja�vmC6d�
|��g�n�<!�	�M����G�}�P�
gKJn�<��B
�b�P���~|*��Dm�<��I�$0��	�����ҵ��q�<)t�̱}� �jbH�N������m�<���F�Q�"(2�SY�\6�f�<1�f�74L��
�N��ܘ�/�`�<9��^(g���0'��",��p5� T�<!Uk�P���{�Kʆ.�½���_O�<���#f�R+�.�7�����FHa�<���G�ꅪynV�� �g�<� ��2q|���O#m��vlf�<��bU�4Kʱ����1��̳C�c�<!�%�q�`!i#�b��!'�E�<�f��
��h��.��py����}�<AFAI�y��,#b%e�xG��n�<�f'��6��!��
'<ͺ7'�j�<��/eO"y�c��Aa,(6��`�<15e] p�Y�c��*1���%�Y�<�A��"�l���W�5�<�#Ra�<IslV�W#��!uFN�D|���m�x�<���q��]c�=�jE#��u�<��Q&u��I�gM�̌k�'Qs�<�g���z|�fi��Vx��� e�<a��Z�d'�\CD�P>.]�� �a�<!����\���߻X�J�3��c�<�B�	�D�"5S��Q6F4>�6�I�<�f�R�I��A�߸��Co�<��O���p���\�����,j�<	���AL�h��k�[Ű�*ŇJh�<)�B"E�y�ՃΒo��U�1�Fd�<��(1Wp��"���^��f�]^�<�HZ?Y��xAgq�mbD��u�!�D�Fc�����&QZv��pE��D�!�$Qx�%���X2%%j�x��ș4�!�ē6p̑�b�'�<ت�m<:�!�� 0���6w"֕і����l��"O)A�H�q�\��ŨR�$ ;c"O���C��.`�`�ԁ=&J"O(��B��N�t����Nf�}�"O,�d�S�z=��!N0x1^�0"O��F�ƫͰd�5�b��t�"O��j��P!\���$O�f�Hs�"O��BJ�23��{�D������"O�\V��!F�:xJ��͗ ����"O>9P�l�+�B�+W�X�)�P"O�!;�+��6�]��u��T� "O2t��#�~~�0e��M��l�u"Oj����M�a�qU�	u�n��"O ����?>� ��员Xc"O.��1�N�	��@P���*7Y� �b"Od!�֣®e��A1*K�s�f��E"O�={F�
V�j���Y�����"O�����:��5"ɟ���"OhhP���Q������>�
]��"Ox��M$ C���DʊX���1"O����R�Feܰ&��*�h�"O�mH�gH 8B��!�Z��"O��KNR�:؛�@B�戨��"O6��W��84�\�)C9�r�"O֔��*ۯ[�l��(\�1���f"O����ˇjDb�PF�DA���A�"Oj< VV�qA"(`���!��0z�"O� H7Y�v��	uW�+���"O��F��K��}[�� 6)q1"OV��_�RV�F� \x�q3�"Oĉ�2�2 ��փ��Qt 5�Q"O�`x��
�@�&�ӄ$�si����"O�,�V�$�4�����*@z,p�E"O�lɅ��4�,�z��2J�q��"O���䂥%q�`c�R6,�Q��"O�p��T�J=��$NҎ}%��C"O8�*���,7n컠M[�ak"�#�"O�x��drbH�PVP0@"OvL�E�ףwM����A�Xܶ�"O8�J���V� �hq,��slT�6"O�Jkڽ\��q!ŋ�$dJ �"O�� 	��I��YĞ�i�a�"O��"O�F#��;��$IN��h"ORP{�l�8F:H�(-"B�j'"O�-��bJ�vd�92��5L1H��"O��5A�WE,T���F*�)�@"O ��D���V��i���5H��i�"O����l�8�F4�F�ÈH��["O�Aa�Րb[�e��
"����"O�h�a����Ƞ	F�&�����"Oʸ��F��(�?�6��A"O^y�WFʽ"*�	�V�X4̺���"OBH����u����h��5"B"OZ�;g��"QE��S�ϑ��n	�"O"l`f���%��n�&wxL�'"O2�2��ۛC^��т�]�?I�5��"O�-h�#T�`h�ŉr�%%F�	�s"OzIh�4%�����D�W���s�"OH@Q�#q�ӣ���8�р��|�<�&�B��:���O��b\v�<��nV��S�K�
%���6�s�<ɥJ7�fl"������t��x�<��)�.���k`@*<�e�[�<Y��?���JT��w-FiX�! V�<� �,�ԝ(!8,��BH�13"O$I�.T� H�9(��4QU�!��"O|����BlXz`����MX#"O�	��҆=[8�b�:��Y�"O<£,��T�q`N1��UP7"O�p����ɐ�� �#-����"O��� �<6���Z"
��""OvJ���?4� �Rm���ecW"O�������N�8��	u�%��"ONuHc�B�t��̟E?� �>��Xδ� ��T��{�1��ȓiR�(�LU,�Ya���~�f,��)u6��g(6��PFO
�T& �ȓ(r�hu�=-�Pء��ƕ(r�<�ȓT5�SRF̚?� ����K�>��ȓlr`7	�M`�� ��"⡇�0.d��AĂz$&m��FM=-���^NE��/�ZW�h�ao�5,����Bq�dȹQ��1�2KS.;p�P�ȓ1��5��*�/0^5��c_�`/&u��)���ҵ��D�J��G�S!�ȓ]�t�c
��\b���ld,�ȓ.K"�*!��%6�dMQ��u|29�ȓ?�����:��QB�L_Bs�`�ȓa�xth���=O̱.�{o≇�db�5#�%!_�"�p�0U�x��GX�C���g� Qb GіL��u��P�E8��Y�s�ʵ�E�Ğ.�
i��K�zTF��w�  ��U�J^��ȓ}6�1A����#T6l�E�X;X	�d�ȓ]CT�@��);|�i�
�=ϞQ��3�~`h�<LI�<c%,G�U7`��pq����"�+k��E���\� ��@��1��K70�a���S<'��U��r'J,Y��P�P܌%R��̷	�X��{��@)�eM�qU��0��	^�ν���D�[j$iE�q��S�%>$�ȓm�@ �����d�=Ah��[h��ȓp	�<ia%�;�hDS�[�|�8�ȓy��lPP�t����-�
��ȓR�,�:�i�Y7,���A�BR���ȓ5R*HY�%>l�D��(3B$��'#��o�g0�aC�&րe��'7(Գp�T�l���TE�"S�x
�'_f!qf ߫n���.̒������y��1l���[���5��<�@j��yB�I�q�V(r������0�C���y��Y0�L�O�� ��M#�W�y�<$ѐ��#H�012����y��Fc
�"@�ϋw�6����ٔ�yB,�
1!���b�j�܁�p��y�,Z&�e�B�\�KЬ�q����yr��+!���b�J�9V_��j���y������@͋OC�)�aY��yB�f�H� �֘>����/؇�y��L�Z�L���L�2�����A��y҉��J�V���E�1� 	pR���y��ܠH<��۲�A�YvN�����y��X�ؤ[0�5#
&%���ߌ�yRE��<��'/�C�z��P���yBF�H=�5���5�����?�y��R�).fX[�1�( (�O��yR��;�6��.��4��`�󭘤�y�M�d		�ɑ�.�n(p3��4�y
� �ɒt�A(¶%�%�	[<��"O���F��>ɀx��꒞3n>d� "O`8���b� RSJ��0e����"O
��US�t�#i�`|QA&"OnI�b�-q8�� (ߦ^NY�"OS�`�,o��I1C���x�)Z%"Ox���S>x����I?�TS�"O��b�F�S��AE� U1�"O>�jU�	T���QgZ�S@e��"O|Ekł�(?w��	A�6>JX`�"O���f
	���iA� &.��Z�"O���ǎT�4���c�,�o�FIs�"O(5;��x�9�J�T��������y�m�q�*`27�[�鸄��yR	�ibL帀�Y�ܰE^:�yB�K�21"q;��.$�$��G#��yB�ȨU�x� ���pH7�U�y�?1�\PRp��
歋���y�f\�T� �'Q�|O�홇-V�yb �i@�)ai�r��x�6i^�y"l��,n�5��,��\��aEh\��y�\��p��ň�)FV]p��ۙ�yn��m<�����D��$H�����y�C��~�	�.�� ���Ɗ�yrE'�Ɂ��Wˢ��TL���yB���Y��լ��N�Lr��]��y�+U�E{� "M5A,�à�&�yR�[j�`g]�L��}����y�ꊰ!n����
X�GABM0����yr��:���A�?Cp!U� �y��\���u�R�U�m�d�];�y�,�1e�t�je��N*~U1g,���y���H=� c�J����V) �y�M&g�X�E�EQ�-P�,�yrj�>zuz���m�A��!�yBi�H�n�x6�Z<lc�AV/�j�<��S�wH�K%l��ZH�2�i�u�<y�.�8� h��*&D+f�n�<�3�ڻn�|P+ �ػ'%�Pp��m�<��1�����9�>��d�<��cKMpj̲�%G<5��Y�-�K�<���<��(2tk"�n�<q�冢F��`���g��P�(�E�<	��Ґ<�(0����깪w'~�<����g9��qTaV6_�|�@B��<�!LO� ���U�(8� �'�{�<���N�]�&@�/�-h��y��#P�<!�iP$yD�A!���pbZr�<�'I�_��5A��Ll���+J�<�g#��
!��r�	ة Li;�cA�<W� o␵@��"B�ɱ��z�<qǌ�,մ����C�D��Xa�<qb,�fYX=��Í�M]�)�w�Z�<icG�[�H��S��c�P�<�p+��<"�rV��N&Pc���E�<�$!"F���8ye~-�6ĊB�<�F�:��[��Ż��lX��f�<1B-R���䢕�ú"���[�(�j�<I�
2I�m�S9lY���o�c�<��.F�-���E�	�LF�M� h�<�6g���A�N��� g�d�<I��i���7#D�3�-M^�<ɢJҔX�t|AAӫR�4QS� TW�<q$ ۴X"p����gM�#��_l�<� XiY���0y󸅋�f�
%�Y"O�t�0� �|$���d�.�l�Q"O�Q�4�}nr��!�I�y�v�Q�"O��iV`�vT�	�tB�a�6�"O@Xs���#Vtz����ۋ����"O&qp���]�,���m�d}j�"O�UP�A����U�?i�}Cp"O�Yp'�L/$0�L����WYB��p"O2�� �o�I5+ /V�	��"Op�rC��s̬�ҫ
�5?@)W"O��͎�c���1Ȇ�67�|2�"O�< E̜�p�J0Sb^�C��p�"O����	 0!x�Xh��	����""O�p�p'�Jf���U.̸] PqsE"O:h�A�(Ͳ�8>�\��>��\E�8s�3k����֯n���I;����b����A
6[{�q�� � l�afָO1B��nL����������8frd���L�n�Y��c���N V�.`�u���rː��ȓ!�`$�1D��Z∴d�ۻ;h��ȓ$,t�1��9�D)Y�K_�Tհ���}5,��W,rW�Yѧ��恄ȓe�I�E_�Q=��Pa*
�'������hO�>ua$[�f��i(UƹP|�b��8D�h�q(	���=�cƕR�ԡfl)D�Aхޘt��ď���$�'D���'�������'h��q#�&D�$c�GC!jYP�3S��d�&d�S�$D���Í/2���xećuO�0�?D��P�ېx�T-z��C�2e���1D�p{oՒ8K�I��_�C���3D�8�uKI.`����5�� "��1D��9�:woF<���HWklbFo5D�����B��$2�Ɇ
7/j��2#.D�� v&@��L(��X�Nf�0w�+D��j\�@obA�C�4 �m�0�,D�@Z���'5H��p�˅o®+ l/D�\Y�K�;��P��
�	D�4��h/D�H8�꛿L����&�I�"HQ"�8D���/ޗ����s�U�}�� 8D�H�׬	s\,p��C]��0 �#D����J�c�a�1��M��,�Q�"D�L2�f�h(j��	�|'i��!<D�hh�C�)X�����@�&�@iq�8D��;ÅA����c�[AЍ��g)D��i&��~mc����(���+D��q$N� I��4`P�n�v��
Ó�~��$�	<ؽs��ϞVk@DK`ꃵ:7!�d؋e:ڍ��/5L_��"��A�X!!��_83�9U�υ4�vAڑ(N&Tx!�ĝb����g(	�	�R���.�!�D�Z���4H��x�d�����-^!��Pw��2E�+�4��5(H��!�d�N�<�9`��̀v��p�<I��'Y��2��a�\�r���R.�S�'�J`�c�����po�I�� s�'ؾ ��.�/DZ� 1�׽H��3�'"��j�A�29*����=��i��'ŰU�%R�Ix��'(�>�+�'5:����|�`��<v*��[�'^��8�ѹ=K��pa��#j�<�b��W��ywW�ZTB�T��`�i����yB��#x]�i�w ��r96��g�:�?��4�O�#>� P 2�A�0�b4���N+x��d�T"O�\X�	8��9ypn��BT&��"O^��W�=��y�@mN1: ��"O�c0!#�h�"셢Mrd��"O(5�D����0�$:fЕqS"Ox4��'ƍn $�jB#_?6�q�P"OjUIe�7Zu�:�dR
o��x� �k����h��R	VqZB�[�h���(D�Pp���A ���$�܆zԚ�:�&D��:U']4{��9�b^�?Q8���?D��ㆨ[/[ i��>u$	�Q�2D������Pn��a����aG0D�\�D.z�T�ʢ��B �)���8D�|Z���%]�.��mV�,{�.8D��9��7~*�š�*@c�4t�V�7D��Kd� o��m�!�]+=uXi���4D�L�q�W�-<��U@��X���C)7�,�	R�O0�� �N+$@ļ��Ú8�|
�'����G�Q
؂5�B�㊌��'9����3c���UG4&R�@�'�� ���)� ��s�	H��`c�'�v�ys	�h*�-qFD��9ܒ��
��y�dS�C���T�Rg�� B�ymٻy_�}�Ā¥Z�����0<�)OʒO�C���*g3�6*݄�i�3"O��	���
OH��C݆8W��P�|��'���ӈθ
�NE�7e�l�H}�
�'��Ј���txԎL�f�K�O�I��h�>)Ó��8�FY�
`�!G�������M����5,n A  �ky��KP��Z�<A )
H��thX���Lc���T?i���S7�4�R�R�K+�@�oҙd&C�	J��� ��5E(��"	\�V
�B�	3lRڝ�S"�0n�yf�My���*�$Y�i2h��^�Q-�E�L"p�!�D�9~>1��GO�kW�B�t�!�Q/q0��B�B��.�5�!��֮~�T��E�ǜ^�<d	�LZ�f���)�'U��p�`�n[v�3�O�e�N���'!Zl���2���P%��c�����'���i��6`���(\�[��(�	�'�j���#�Sl��[��T�4��I>ш��)=@��ӌ�z��x['�S !�dQ�"�\�0c���*��C08r!���%!��E����&w�A����2n>!�B�I8�9��E�HqB�
���!�	,kq�H���&Y��BA�|�!���W�f�Yҫ�Am�s����
i!��{�e��A��.�0��bO«M!����$ɰ�O��'R��/H!�	%d�xUr0��Q���K��!��=��`J9,�2Pď?�!��P7,zp��搏6*�xC��o�!�"X���gLL(@�h���^�!�DJ�b��0�S�҃vk��{�:�!򄑍>A�(��O#D�f�jℐ8 �!��3
/L���d��Q�u(!��ȟq|��M�v�~D���!!���<������k�v\XՅ+o�!�ђ:N�G��=t���G¦hU!��� 99	c�`g���DߎM!�D[�y�XXdl��JJ8m��`� P!��4�r����I�^F��ꦥ�� $!��H��aC$����ԃ!�� |-CF��V��#���#�	K�"O̠ڀn�"Qs"�c�`T 9�g"O�di�/��(�F,0����8�s"OXكq�E�fi� H��M�Є!�#"Op{Ȇ{*�B�h��ik���f"O� ��߆0%0�Ф��V�$ �"O�:Qй(Jd����+.d��x�"O��+-���z=�6��dÎL�"O�͋��9V|\ZaEP���Pf"O��c�\I�!��$�(���s"O��q�H��[�f̥w�.T�f"Oƥc� ��}r�AJ�J:E���"O����-O�\4��r�yM�
�"O����-�Xj<K�
R�q(�"O$��wA 51b�
E>;7�<��"Ox �*��tM��� L�_,�僴"O`�3�Ò=4�#��"&~�I�"Op<���j��� ˔,L�*�"O��sD��|<��2H��A��"O�r�f���·�N����"O�����#Mt��e�F�( [C"Oi	�&�{�pQ�c�	z���P"O�r�+k�`,�c\�7�A�"OL%�C��S䴍�@"���V1Y2"O�d����V
��L%Q��@�#"O��K%C���ڀ�bnD�#�(-��"Ol8q��^7H��b�\I�肠"O-����	��$��lS�@D��[""O>��VbY�~!!�������S"OV�X!�ђ���
�X#J��	c"O�k��S8����#S�S�b<��"Ot<��E�#Y�.�h�E�L4�U"O�0q���sK.�r#��$|<���"O��@�]�%c�� ă�;y�٠�"O�1�v�\��X��CY�K `p9�"O�� ��Kf�0���� F�ԍ�4"O������ vMl��4*��T��@��"O���됑 [z���iD�i0R"OR��O��NR܈��O*t�"}j4"O$@c��m�5��\�i�6��"OJaID��25t�H�'�x�`�"O���0N��= ��(�b<�"O��kƍ	�y	�Q�`�%j�Z�X5"O
��ğ� xk�K�B)���"O�TJǎ�q���7�'L���"O$�B��mzZ�S��k�&��t"Ot���!/�)a�i�)w��A"O*`���R�9&,X�DI
<e�Eib"OF�q/I>>�B�ۖF��wߤ���"O6�B�nO�e�ڙb��3%v *"OB�3�!G,Αx⢇0D@�ih�"O�pK�b�2l��i�SH��}N�B!"O�Ѹ�G̹R�m��HC�	���Ѣ"O�L@WĖ�0�I���@"v�F�:�"OZ�C�(V)Q}�p���;m�,�"O�R�ƛ�`ց�B�_+dO
��R"O 1s��c��"�2"rh�D"O�tJEH�'TB2���ۦ.��$Q�"Oh�[�@�;�lС�T�S�Yz�"O8�1��ߥi�r�	)�5a�Dx8t"OL��'�؞k�l��P֫\�&��#"O.܉�lr��!�$u#�"OL���ጕ@��`�U�۔F�ݛg"O��2䢘�w����熇a�De0�"O� �8����%��tr4eX�@X�ig"O8�e�(�68Ze�P[����"O ��ƃ������	fQ�5aE"O�m{��-~W>��v��d��My�"O|ZV+��)48���F���,���"OXqF�E
q+�>�A�p"OԨc���/Y+��x'��DJi��"O�e���S�o
h�;�^5�E	d"O�%�b� ����e����&"O $A"H��mA�^M
�T"O����J��0�������b+��e"O1G()-����N:D��*2"O�ܹ�k�{
&,kR�M�DGX�P�"ON$)��~�:sK�K6���U"O��J�%�r�"R�I�BF��S�"O�,��H�!XB��E�7>����"O���b"H�O�q�ĤF�c��¥"O��'C6xH��"䄩}U�"O��0�r�qU�ԉ{��䂲"O�7��("�ؘ�@Y���@r�"O�����Ga�H��$~�z��a"O�� �*�� �lh������4"O��a6��[Z4����q��m�$"O�p�cҬљ�>gd��"O,��1��\��o�� T���u"O ���B�^x����ZGNdhG"O���d�؎dqh�a�#Q ��Y[�"O¬	��ʡ8�x"�Χ� 	k"O�x��N#��h�"O��6��P"O� {t-��Ba�S��+w�I��"OV��7'�w,��gKƲ�ZX�"OԼk��;[.��r#
� n��a+�"OX�;GA[�#�����R�7eڥC"O��t�ČV6q釂��PI�-��"O@QB�)rVp�P��L�L�Tt�2"O>����${�$U�E�lö`w"O���c�
OT�z�%�*\���Q�"O��Y��U�F��K�$�����4D���@�a��-�6�KEe �su�3D��rF�9n��(��H6�5�ת1D�DcCEkh�v
 @9���M1D��ن���4VF��p� j�U�ub4D�(�ʓ��쳁돥7�� �cj3D����e˘F�|u��X>ɬ�B0D�d�!X&>�@��%��#~�9��0D���]�"�(mY')��F�)D��8�Oگ9G
5�&D�܂֪3D�L#ʰT}ԙ�%�|�� �1D��Bc�"m�TQi�O��%�4�D;D��Z���S��5����6��Ag�:D��k��b�Z��ӓ��1Y*>D�#�L�),}hx��OQ�&"���
;D�|J�N��F��9a����<��m5D��qt!������S	%%4qf�-D��jգ,E��)e��WZСӒ-+D�ĐC�
��u
���"n)D�x �!,�8��d�h�I�Ԧ2D��hn�?��$�&��.YYB�p"3D�2���Lf�a�aQ��Vdɀ%D�@��g�7rҥi�ʄ;	v�)��$D��T�B"Ew���Fǭf���uG#D�0���ʬr7n���4!��4���"D��J5�CSN���+x��DB��+D�,�w@�1��m��CD8�ĸ�..D�� �t��oɐ{�*1@&R�R�1c"OH��C�[�*�|�k�D�V�"��"OX��0� �1)r,�u�¾N�ZuP"O��6�3H��L�+��i�p�r�"O�	��W($h�u����,Y��"On��+K!O6�(��O<�<�S$"O�reGZY90��4ǁ7d�Z�"O.=ʣ�A"r�����E�95�\8s"O`|��Z��N�e��5��A�"O&)QC	��6ц$����;��P�"O\�q�f�J��x�C*ց�r|��"O�2���_�E�e��67��`@5"O<d���	#K�Ѡ���1\��\��"O2�!�$S�k���" X�BL��!��¢|�N��$� gA���*H	!�D�2���BS�WA�Ȃ��̦�Py��2,T1�"��wP���V%DN�<1�ED���:G-�!ӂGUf�<�B��Pj�ݳ �J+�Y���`�<q%�&"�,��Rk'z&��!��Tr�<��*�nePs�P&8�8A-�o�<YS��
I�^��à#Q��-+��g�<�aK�mv��p!nҜ/(�	[�Ee�<Q2暑*l0X�J�Y�D@��_�<��'������5-Ux��)Y�À^�<�D$�u9 \�"σ	t�`A�n�@�<�Q�5+i��bU�8����y�<��ڿ}	*�;g�]FuxE8��}�<aE�&>��� �k�H��Al�a�`'�|��Cx��e���_�!�wB!D�;��J�B^��(��>���gK?D�dс�=��yb��]�/6�p2">D��)�FN�S���ң&Z�p���B)D��`�" �`z�M�r�V������(D��;�A�C��2�f�OP�8j�!&D���6N�d�b���hN6>��i�c$D��Č
�yl� ��H�W.5R��'D���E��b;Ƒ��d��[��dR�@'D�(`'T�xf�M���ȜF�4�X�&:D��r���'m@0t�	��pW�7D�pz��	F�(I�'K�#AX"��W	4D��	'ոeUpp��ìt,Ca�3D��C�ޔ`��4�@1�Yv��Oh<�b������������y�F�'{����D�.# <���W��yra�"���'A	-�q��ș�y��.���VnG	9D���R�3�y��=c�NI�vb�24��ІD�=�y´l#����@*n�Ŋ��U�0?�(OzЈW(Z)�x9C�U�^@V����'e�OuQ2�EL��U�����c4Z�A�"ObPsR��
.�؄1���r���"Ov��`M
@���� H|TȰ�"O�ESG�PQ�4y�֭&_���ȑ"O�9��Jбfд�I��o!u�@a�!�$ψh!�� ��,�J!��'V�!�då,��Q��W?H�TP�L�E�!�D�@�����./���BMy!���'^v�ڀ+��a��=�P!ģYp�$5�Ol�Q�����`�h�uf��{�"O����� ���FҐS�hH�"O�Z�� ���Z�IVG�q�"O�ҕ�"�U���؉"4���GO>�$�>@g�9!�;.U��-���'�ў� p�jA�';E:�c$@�y��wO��W#[6�"�A�5����$GX4�!��\*s��	fl!�hB䔲�!�h{SLԓ�	װX��^/?�!�D��8'b\2��6i���"��\�!�S�z����""��� ��`�!��R+N����J�W��y�`٢	�!��4[$�Y��˿x�j���L�	k!�ΚD"=₏߯?�x�)u�ՖT�!��'Y���*��� �0�<7[!�H{���%	ЈM�*˸x<!��" t�
s�)�b◩�!!�Q�^�\ɨ��ٮ;�ȑ1q)C<\4!�>��tۇ�B�
0������3�J���S�O$2�@?A�<�zw��8uz ��C3�y��1@d�1"�/7_�rd���y�U,Q*��	�e�Na�e��yBb@P.9��bA�n�(!� ��x�<���GK �20d5��)x�Nl�<��Ku��-��j�3Q�~��"EE\�<a�Æea*����O-<z�8xAk�^�<�4����x�@$bt�0-�[�<�E�!.ي @ cT!M*�x��EOT�<�V�w�Z H7��*��;�.�i�<���<��M�a×p�v�2eCTc�<y� �q�� J��A8Iy(�pc&�`�<�#�B*L�Bq�L��X���_�<��
�y^H�g��ID�h`��OF�<�Q/#h�����#��(q�B�<�&ĶH2���D� ��`���<��@�dP[�F�^k�б0��8Tr�ȓ9�@�(6��c��`�E�i��ȓ\q`�ke
��:��q��42TD$�ȓ��@i�NŻJ�h���R�Ed�!��lsJ�1��Y�3�ެj1ϗoU��ȓiIN,1TIРx*虇ኩY,��Ju�ku��{پty���!�h��<������O��`P�� ����e�@[Z��	�'�T�9�凂9Q8\YpO�.={^��	�'�$�S�h!@�<���'�~x��'g���w���C#(�b�ɯ+kX��'�.���	F�!r�h�O�:*4Z�C
�'_:��T�:f8M��/� �>�)
�'����+=�MȄE�N�!�y�S��G�C�UqnD(B���F��XcGJ�/�y"�#R��r�lö9�
��6O��PyB#�1sd�x�GL�#~�|r1�h�<	�"�U��p����[38)Z �O<9�r�&�� �1X��4@�vK�l�ȓw���Z1ˬd4� 0٦��ȓnl`D�C�G�'�0|8�h_}P�p�<!��?���� :� R���8F����K�D !�X�/��@�v�Y������Ƀd!�P+%�ᐠ�11��	�i�,K�!��%����GT9nJل�=!����
������,�C��B!�$?R|���S).ݒ�x� �6M�$"�Oxh2���%B6:%qT�
��q�2"O�2 V�PL� �G-�"R��)r�"O�M!��X���wX6,�>�� "OP�6/�Dj�c b�����"OJ	�� [�!�j�á�@=o����"O�YyB��)<yv��捝����4�34����C��`�����!aW�t*��:Of�=� Ё*6��$/�l�� gI�0�T)��IYx�d����o�p-	p��1A���8��*D�X�6�K0�� BA�}���F$D��г�3rP 9Ф��*�1�!D��S��v�r�b�#H�$H��R� D�l��O�Cz�2m�^ʬ�c!�??!��$,���o+T̩�	NL�0 m��N�B�%�|�{3+"�x����"}BB�I�i&*���b�jF�YMU>�6B�	%�U)��� e�*�j�j� &4B� a-�[�A��9i��� oC�@C�&WxX�y]Ep��g�țY�P��'�l��F˝(m��1@�_? U��'�N-���"��ڂK@/S�Y��'Hn� ��֖Q��٢�B~Ј��y��)�63��R���$
j(特��B��{u�	^c�.x"�K�؀C�I�,
��p(F:��O40�jC�	 ���B�MEJ�ᐆB�0*�>C�ɪ?�X{U�	74F	��	K�[��B�z^Cs��5m>��*ǆ~n�B��$���&�\�)��pCX"jw���hO>A�&Eֹ8�u��I̊P Z=ac�*D���vH�(Hix���IW,2،�[�G)D��{��������	�(��bG=D����M�s~D������`'D�hsŎ$f�6t��*Νb⤝�3I0D� ��
yЭ0 �rI���A++D�ܸ�(ڔ$�8j���J�9E�*D�Ԁfi�.&>�� B��
!��+D�,(t���9z!&:"* �*ac*D�И �W����"BL�]̨P�&D�0�CFN�Paj��U�(Hpb�
$D�p�t&ցa�(|��Ƈ8U�v=�! %D�<S�V�s��'�a�
Dr��$D��0d*N(	�Zp���1��5*4+#�I[���� ��/Tr�3L� �څs%�-D�S��Q���JFAH�-`���(+D�Pk!!P!)Jhb僤5��(ah3D����׹]�q)�>b[�E#�h1D���X�Ψ��"��_��\
6�Р�yB��s�'��@oZ�Z��H��ƗS8�e+�'f| �D�6n0A9T65�.���':6)�#O���ܰ��O1�ҹ�'w�9�QJԣY]$[3D�2O�@��'�`T7Oؚ+�lUHcM�$xi���'���+�9"=��FE�>� H�'�	���cv�3�
ʱ~]J�3�����XP�S�c�
���j9=�Τ��#� Y���4fŚqR�̬F���u�V�(��N�q��؈���'|I�%�ȓ4a�h�g���*�`�x�/�8I�-�ȓq�V�`�3ih (/H�<R�ȓe�d���9<~xj���,Zt�u���@`�3B��-
��3�p�ȓq#Ę��%��D������W�T����ȓ&��k�Kcag=�����y��@�ץ^+7�"�!%F��d_�`��/���� l�
�YB���t$��B�.3@�$�V ��J�!VB�I��ة��W67ĸ�AjNvRB�I��Bh0p[��v%���d�X��D,��_���-Ir��T3+!��1t�99'H�f쑚��"���F�� ��8�Ϝ�R��Qcㅔ�i�2���"O��J4+�/�=����6ec&(Z"O=	�/�]��|J""�^�@a�"O��3���a��,�75��c"OnY�!��xp�)yS((*�
"O�d�5
�4+U����H\�f���"OJp�������{��F#o��A�q"Ol���\�g���mT�B�M!`"O�e �2b.��&���K�B�[�"Oި�F�Ь0ɰAC�kE,lZ(��"O>� �ѰC��l�h�:(LxSe"O�<�&j� PY6�Å���/o�-{�"Oڍ���>z��dra�K5hn���"O�0!5e�@>��0∖q`��ǡ+����"|�O�ĸ�F� nn�����,o`��'�6�z�-E�nmi�Ǐ%��A�',���#��Q���J�ʛr;Z�	�'�lt������K�c����	�' P���Pb���EPG��0�'���I��
�q��a��
*�yNۣ*p��H�]�ޱ:�l��y��B�"j2= �*ӥa��l��͓�y2�O�\/�u���H;_��x��@4�y2�tY��0�M׃U�vѩ+_��y�^R���NI:HS�t�ťG)�y�_�?5�2џl�$ᴅ�Xў"~�-I��D���17p�2�$t���ȓ`�4K��N5g��a�v�f�bi���l�'Z����ʀ�a B�W�*�X�'ހL�Uo�dq�lԠ,��'�D=R !ͫ¼}�B��
�iA�'�Pzg�Q�
Q��H��p�J
�'���VXN�i��[+}c�U@�'W��K:~��:S�	��nt���Ƽ�yRݻ#�b59�	�M�\�#����yRc�v\��@(�н⅊Ò�yR��;�XX�K(�Nՙ��L��y"��;0FL���AJ�5%ʘ��AVv�<��h�(��m�Ҭc)r���W�<!WL��i`f$��%��\ �B�Q�<�"Q$��{7NY�=ᘼ���PL�<9���<�L ,��%�pZ�N�<��9)�L�@%XAl��#�VC�<!�-ϧ8$�k�/ŋzZm�#��~�<9ǯ�!b�R��Um_�s��X��w�<p*��%(򰠡!	x����G&DY�<I�n��%��`A
��sF�Q�<��a�#6R.���?(�r���`�Q�<���e���k��l�P�[�)P~��)§b��}H�
3<��ݺ�U�#"�ȓb�B�j���j�����z���ȓ:_� ���A�C�2Q�EJ�8��ȓKQ$�b�O�P5XL1)�#wz���za��NY8gp�$Y��,���ӏ��s�|�)�F�R��vɞ�|�S2D� X$��^y�D򒋅/ 6\�@5�0D�ԡ�@��+�Τ����A"��Z�.D���e [0y����F�>�V����>D��sR�
r�p��$e>��v;D�
U���m����~�۱�<D��Z�Ӄa�1�'�M�WߜT��;D�<��� �6��){H2%(L�7�7D��qBɠ[�V�r�H7n*8j� 4D�@ C$>�ժ�kơUP�=D�� lͨ ݧ{'�٨%m:��2"O0= ԊT��D�Q���u�m��"O}�7�H���Z6e�c�|���"O���6��6�lA�!e�="���
Ō+�S��y�Ȟ�@�Sh����A��_��y���lhlx*#*D�4!4xh����y2(&8�S4؞��v,��y�ǈ$mP�a��`�%	o����K��y2eL���A�(Kz53.X(�y�A_/��qIRI�<�����Й�y�
:�q���^�C-F:V5ў"~�ENRlc U�8�Z�su��M/>������x��w/��ҩ4����"�ܤRm߉i b�2*��`&��ȓL����  �s~�=�ao�kW&�ȓ�8�(_�
��a"Ҋ<����ȓO��툁`�&s���#ݡB6�d����0R��>��M�7�Z�u�4��ȓw�ص�̕�0s�X���@7wR.X�ȓ���1+\o�XYң��\{xx���&�`�`\�G�|� ���1�\�ȓ.�x!z�A�7;�*iw#��fQ�ȓ7,�3�#�0Ĩb}d��ȓs�`�1��7(�1т ^.2���ȓE%扊a�G�]ȅezk �ȓe�8��֡Q�xE�"� o��I�ȓ`㲨hP�"(�����?a�|��!���%Ȅ���K3/ �4��Ʉȓ�r�H�/�!�$��td��N�ȓO&�̛6�U�Z��i�� ��ȓ3���䆕 �|���$8�֡�ȓ[��(�����<�!	�vSԕ�ȓbǔ�1v	F�F��Mj��-�ȓ�T�#AO��!��$��}�r!��?,y�͈4,������&9��n$ӗ/ֶ�L�Ӆn��h�!��+ �te�Ѫ�0�[ƀ$��@Z�<	am�)��sW��Oq:��%N�<��h�Z����phnAJ��_�<iUȪ:X�(����9Z�Jw�<�%Ɗ����� IV	A~L#�e�|�<���B�yu�KC�W)U����,�t�<�0L	�^�4�`X�fZ�<*�mi�<���'\��5��uL) ��b�<��M��6�Z���i ��C�ɊV��H�`cɅ �cU!>|IJB䉣"�N�!.�1��l��3j50B䉋i5�%3To��U��ȺQ�� 	B�I�L���s��ٖ"���bF���C��1/��p&M�4��Hp�m�*,~�B�	�Oh�����\�a��}��b�*N�B䉝mXГ@�Υ�ґ��iԙY+�B�ɼ ��p���I���2�`Sfe�C䉂MD����Δ$����BS<��C�I�d#��`HB�,)$VXB�C�	"��Ѓ4.B��z� e/P�l,�C�I�s)�a"زb����է�Qz�C�	� �l���M��`�*O)z��C�I��KÃI�b��T1�)ȸ y�B�	�f�$���cqhl��X�ܸB�I1t"�c;+d 2$�U:hC�	�("���n�_gT�p-�0eB����!f��&�|,h�ϘoBB�	-u����N$ �Ta�F�/n� B�)�  Ha@���h��wiH�u�@��P"O6Ƀ��ǆ=�z���5N��)H0"OzݻV"��[+<,ˡ�j� ٸ"O��%��aMB\�F�F��a�"O �$��6�L�Ԇ	�b��4ڃ����II����s��t�+��kA(��H1D�L�`��z���
ͣ��k�1D��:7 P�v3�]�G���ܰsJ1D����$Oe��j��nʠۃ�/D���"`I�oi���KH)�diS��.D�L�%��8�8A�6�J�V���9B�+D�XF�īw��L�F�〈�k,?i(O��$ҲQPhJ₋�;I6���l	�t�!�+�2 �N�89p�8#��&W�!�DV�4���A��,T8��Q	��x�!�d�
,Ӓ,��j�5G&��ZUG)X�!�$�	�,�sm��f���Qq`u�!�� ;1�$A� �H�	�
X�OD�#�!��%F?t���F�Yk4�����/�1O����)����ń��]��KD��){�!��<&���T�����{��E$+�!�$��8r�l�7����"�(�KH�!�D�m�̩���4l�P�1l	�x�!�$\�2`�� *�	O�1���W�!�D��@���B�]DA�U�k�?W�!��BR���,��#���s)�.=l!�D�Rq���5�[1W8���!HN��!�H#1�}���P<	C	wGP�*�!���h�8"-��t�%�7�S6e!��ZcZ0�[�e�='����MM$u!���}�d!x��O�a�+݂@i!�DE8���AL� w	�Ũ�^6!�$Q��h���o�L�5J�;/�!�dl�M�S�
�%&T���I&�!�݄�+.��=��E�:?3��ȓC}.�4��/�����띸.�R���X�ɪW=�+V�<*����DӦG{��9O�  sIR�b#nQ�e$[�:��ɣ"O�I 4,��*�qc��C�z��"O����E�j~^����U�:�"OdP
��3/� �(�b�15dɂ"O�u#�-K	Z�R�ݏD�슗"O��xq��5Am PӅG�� ��&�'��'nf�7�u�
�����}���j	�'2j�څ��/jq(y���{�ą	�'Ԋ��0���k���i� ��:�R�'���c�W�B��[WO��uAl4�
�'��'mA��]���K�Y�8d��'B�A��f��<�B��;Pm^d��'e�Yx,��0H3j��w$�)��'4�M�` Ƕ�:h��.� 瀝���)��<	RB�X��<����82s(��UQ�<I ���25.�1��5zId����v�<�p��^�D�PU�ͰD;�iq �p�<)w�ުY���0��B�B���0&a\E�<�1���>9�S/.�6a��~�<�a�@7_�m�a�ω;���Y�+�w�<����~���!-
N�,	BG�p�<!��-@�h����VB+��)�!�*p�,��AL�^�{%�B�!�$ܭj��93�M8l��{�_�s�!��}ځ)uK���JBc�n�!�dK�3r�H�1��/J��q��^P!�=~0*5S�#]$h̀�S%�R�)P!�� Ls����vi�r͕8;�P9O4�=E�4(�vJ>�A���b@�X�!(�y��&Y��8��Ȣ[�T��' �=�yB"3BbV �M]�\��B!�y2�A�p5�y��5(�	 rIV��y҄:$ޮ������́A`Q>�y�*f�v���gBw�@bЗ�y���x!���b���w��\CIî�yR���Q��l{��'��<�yB��6MN�M�@�`�l �&��y�"��@(J�!+C�5�yr�0r̑���k�daɢL��y���_rR����h��L)C��y2�9fD媂ge���aO���y��Ⱥ+ 4��5��c��˗�ͪ�y�GM�!p⸰eJ�#W�^xѧ#��yB�:EB���' R���gɛ
�y�a78�����D�бQl���y��	��ܹ�A�<��t�W�ٺ�y�E�*{B�듶/
mzp@]-�y�×�DM�������1D�5[A@��O&���͝�0XD�%�J�X�˓��K�<y�NR"1K`�B��c��˔�F���?��̉�	�X�B�Q�>0t�b�
�~�<aRf����%HJ�A�R}:�a�<a�i�|�jA'.��a��%����H�<A�dܶI�zI����%~� "V}�<�_"r0�]�`�M<U�����s�<	Al�
YZ��W#6Q�Α�g/���hO?�!."ٳ3�H=U�4��0aK$92ZC��b3,��r7YgZ�y�lH?>N@��$ �$.�P+�.�1+�� P@�%M�Ņȓ	�x)�A�6
wX#օ۟S�r��Q�B(���3!��B�
M֩�ȓ٘�Pg��%G�$�2���X����?�5�ӽi:���.ma�x"t�-��x�����6&�D�E�U�3&�,��'8����5�0�c�-�-�̴K�'u0M��!�W	�`X(����'�DXQ��L�!��8K�Lt�b���'v$��a�V��Zѥ��N��'��*Fg�7D4��@�Ē �l3�'W(�9bc����I���;�H�'$|�P��5��A�>��2�'xƐ�ѡG�u���J���&����'p�e��IO@B8��NJ$����'��yi�M�sp"T�� �+��qq
�'y���J�f�P��̾-�:���'��aa0���-g�͈Ri�q�j�X�'��p��l͕K�<�B׉ت@��u��':��F��Y��=��lК<���ȓhjr��VEU�gJ�
f�N�i ��ȓO����cY�� ���zT��ȓ-�NTcF��C�B����`Ɇȓs�+�H���
�R�(#j�`Ȇ�E��Ě�b�8~G�Q��ӜK����g�M��W�:����fo�12�|�ȓn�<\��[�!��=(��5$Q ��ȓLB��s�["KPL�V�C-HC�݄�{�F� �lr:�c��\��ՄȓA2���`-��UDp��ܦg��ȓa[������m�n�G��&gi2Q�ȓ�� 9ì҃"mP�z��>�6%����?�  �rC (����l�9AP�H�<� �3d���DX��e��]VD�y"O�@R���Yפt��
�=G���"OeB�.�1j�l�'M�/Wt��"O����S)Y���[��S�a�@��"OqC
���]��.��s D�"O�-�0NY�>0���P%Vm΀�"O�8�n͚�<(�c	X[B�("OdՒaCm4�����Mŉ�"O���3%��c��܊�g�+77����"O�A��a���`m���<7+D4y�"O�m+��-�Ġ�hӌu�v)��"O�b�/F�b��A q�ϲ.�@{T"O�2O�ሰPƇ@	d~�1��"OrH��D/�2�A%���|��P�"O�A�+�0iƲ��壖m���"O>U��a�\a$�� LU�+Z�$"O�ã�LQ
,B2D�D��@U"O�����ܒ^�9+���1>����"O�z#Q)���KSC@�w��T"OL����|N�S!�}]R��r"O�L{#��2�d=Zw�+)�"�8�"O65z�N�C� k�L[�D�"O
�)�"Tur���Vȱ�"Ob�(�B�)r܌B	�V����v"OF-C��X�ŢU���if��Q"O��@�K%TX`�i��K�P�"O��Hg��}\�,�B(�>.<�J"O�H�ק\|���6�A+C�Ӵ"ONU�o��D�B4ۓ˚!�C4"O\xP%�X̒H���� ܍!$�';��'��I�)�x`� C��(q�%��7l�C�Ɂ[�,10t�ПB�>$Bc��fQNC�I�]������Z�4����vC�	(%�&p��⃂0��zv��+�VC�ɕbV%%-�)uN���� �cNC䉁��\��Vd/ ���4�4C��!rd���ǌ�*�.�)u���<J���Ļ<�-O@�y����^���X֏˛O���V"O�S�@'-��aJ�/��\�s"O���t���\񈗀']�4���"O  �ˏ&^Z�J�N�V)FqY�"O�x�E��B����k�O��y�"O�Ёb۩��8�w��-
|�	�"O�A@��&unA:"��n)��3��'�P�x
�K�9�$����Sj Ěg&D�T��3q��	����z�� ���$D�hR�'��p����_�T{��0��#D� �	 "_X��'?S��� D�L�� K8�tp2G�M
/sD8F�:D�Hx��X2�DY B�*i(�I�Ab4D�<p&gZ��%�ծ��))&�jo!�d�
�VM��	ݐ0�xPJ�j!��JX���蝆�^����ηQK!��n��A��LS��]�C���I&!�˙Z�ʹ�2�	�u�����"s!�ʅaw�M��"Y�i�N�����j�!�DƓ+��	�`B.�& :E���!�;<<�[�!y�Y0�dƝ�!�˰?^E`�Jg���b�1O���&AɈE�AKU�}f��qc`߄L*!�$�xZPhC��4Ú0fDϻ=�!�X�U��%�0:�����^�#�!򤗯Ffi����`�̙)��S
f!��ܼe���	��%t|�!E=f�!�� ��A�-�`��4gҎ	��Pb"O>t9����0h-�'[���w�D4|Ol���b�3`���z2����B"O�a�ъס�x���B�q�X�Q"OD�;��ǑR�9`dc�*숩&"OVI��ada#��v�B��p�c�!�dY)��T�t�ѿXU������z!��K��C�cӠ-Xa�FΏ�e!�$F�j�lK��r�v�����m6!�˪,�4[vCL�DQ0��ġ6!�d��,nD�!���l1���_�!��	�B�@c:rp����	R`!�nX~A�O�>���!�,Z�H!�Ę�J'21���U�#l2x���q�!��G�� \���R�Gj*X��@!���E 4���	�G��'h۰!��\$#	a��I]�z�{qF�?I�!�dG�>�����#Z�b6pJ�E@�5�!�d�'=�c�R�U�����J�!�D��M�܅�C	0�t�k���8#!��,^@�plm�8q{v��-r!�䀭(�~��j�+}�(SƍK�GY!�\�TK���:S������$P!�
�-���S&��",⒙��	�	;7!�dK�����4!�Ɇ� ��;�!��Y��H���S�2ؙ���aR!��,i��9´��>g���j�Kh!�D^
[�
����^6w��B*4l^!��\�\yt���l�2ch��[Ԣܒ(�!��O_�0����0oS4�#R��K�!��ܘ6j~�J7B�-9��W�T9%!�ރ	�b,
1��	W@�
aI��y�!�d�<JƔ�i�փ;ؠ4�ShK�z�!��A����5A�Z���(~�!��;̒����? ��0��I�?�!�Ċ�5l�0�mP"2��� &H�n�!�$��y��A1���:��`�FU�?�!�D"l���JP.s���ԣ@�Cn!�VN��6kĲ{
L��c �JO!�䛌x�T���P�Y��<����!�!����IY��5�XŨe�V�!�[7��(��L�^��(��ރS�!���0�l�r#ڿ)���L�<�!�[�Z��ę�(X�{�6h�F�K�J!��]m)� �R��r;��Ϟf,!��7��(*2%�%.&إ*�D�S'!�Oi_T�B�x����6F!�ٔS��;����K�B���5�p���Z�)�B�z��$/wtŇ��ʹ�����9��9�v捈*�ƈ��j�L�ˇ+O�ڜ��TG6�`�ȓ#�p։5�D�KM�b��مȓBD����_�[�z�ʓ(�
��ȓ$hL)K*�QK��傂/Ff�ȓ�xhP�mX���GI��ȓ68�fQ�q�8j��$ȺP��r�R��fO�}r��9wP'|хȓMq�=����Bt��KT��Ĥ��~V�0pJ��rn@�N�R�����Lgٛ��I(>LT�B �%T;久ȓD�Y�� �m�cI�s=��ȓN��t��l�I�R��ȓk�`ĂSN��i���@!3�����^����B,H���4�4&Da��S�? x0y�Kȉq����4���A�ڸ�s"OV���U"]�@D	V�L(mqb�p"O����i�G��H+t�Țm~�Z�"O�У���a����^/z�i�"O��!r ϱ>Y^S���;��9K�"O8 � ��I��c��7S��t��"O8Ђ�����B���k��u"O��H(T(a甡�KS0�h�c"O��s�I�H���KНz��X�#�)D�R�L��И�e�q��S��'D��0E�� 2\2q�%g��"��(�a$D�X��F�^z�	�B��-j1Ȍ;D�.D�T8���H  sKn`�H���,D� Ʌ+x�.H���E�R@�qj�/D�lyW�ӶJ�V���F�f�vL��g1D��X���,�I���C@J���5�3D�����A<�1�cǛ�x5D\p!4D�D�a�ݕ�|� ���*1��3D� ���&�Bg��}�䉐r�<D�HЧ&3p�8x�ზI��k��/D����M\dm�1ˁ�46�� ��7D�D�ɀ]p2�"@B�u؀RA�5D�pH��+>Þ�+r+CX�h���/3D�p;F�]�{>���H�?1�,]P4#7D���Oڀ7d.@�)D'z��bc5D���F	Y���2@�>]� ��&1D�ȫ%��q��H���7}�X�M;D��Ԡ�꼈4��	�%�F�\�!�D�?pT��j��&YzW)��M�!�$6	�dj�g\eP��J��u[!�$D��� %�"&�l�9�iU-s4!�$��KЂ8@B�~|��f"�T/!�$��v���T��+jIZ�NNL!��վJ�b��1��C;��*f`U�@&!��$/t���?@G�uɤ�H�C!�d��z�\��ِZ4U�t_��!�d��M�Dr�,���	�W�5�!�o)���ނ>;��95��L,H0
�'2Q��jҲJ��1�,��
�� 3	�'�a8l�as�QKdc0~k�l�	�'S0y���=:�*D+�z�C	�'��� ��/G����ٌ �x�k�'�^�!�h��W���P�� }�j�@�'f��+�S"\TRU#t��I��'Tb�I��� iyƀaW��e��P�'�`4��N<������ZLF��'�Az������q�aFA*K�T*�'�x(���M��d��fH<E�<��'m֭p�j�o�� �叚h��Q�
�'Yn8�.��n��6L�V�� �'�8����,L|�1�P1x ���'��� Х)v���#��hLd�r
�'( cZw�0�� ��eYz�s	�'����g�@X�keO�6\}|���'��܀�,`I�|I��'�"��'����/��f��PV��~؊�q�'@�ڲ,�=BT�9��g>x	�'�<ܨEE&�>�E��/pڨj�'\�1F�ϺS3r�ȵ��.팽�'�� �)�г�#w% �'wf�p���9qnJkB��%`���H�'��z�@�	��"��F����	�'$$c��^�h�a��ǔ0z\���'Ζm"�̗��I�3rI��F�<�  H;1)
���Q�����ʤ�q"O�3�P7� 1����V�b�"O29ӵ�ɑE�~����,b{J\Y�"O���l܄5��	He� jBhɦ"O�eہ�1[��X��Ϗ�r���"O�@ �B�R����.V9T��{�"O=b6��3{��H���|D��I�"O@�P�� $$���F.�0D�A�C"O&$�V��'[V&`qD����r�"OxA� �A���M��ok��c�*O:�B�O�*t`Ibた<8���'�T���!eB����e׻7�z���'���dmՖQ�ܩ
BC�-r��
�'$ m �iY�t��q�J0 �s
�'i�x���NMАiХ�Q�F�Xh��'�D$�� ØOSڐ1`M��A*V���'�~�W�����kwH7ew�H�'���b�	�&J������+��5�'�l����Q�4_�\V揧a�P�'it +v`�,N���nB�:�֩��'2��YՌH�rXV	9��C�2/� �'������y�9Jg��@�� 
�'���J�ʓ�c6�U�8+�K	�'��prǓ�R*Т�"�@:�Dk�'��R&I�P�+r*�Af�TB�'�P���ˑ��S@-��M5`�'�z)S��NG>!h��AN\l�q�'�HӇ�2~ը�+�GE�3�'�y�CĐau�}��k
�:� |�	�'�xQ@�ɞ=:���8&/E�8T�k	�'��Q�MY0%ݰ����,z \tk�'uV\�AJ�- �E��CJ�p�A�
�'�t%!&�G�y�
���H���"�'�V���D��J}{�덳7RL��'��<c��M(ܭ��N.'yn�'������0mH�P�ÉT cb�`�'�
4�����d�d�(ć�l�s�'ML�x"EW�E-��qs��=�~H��'ː��q-I�%(�L�1j�:|*� �'�F�%k��p����hq�j
�'$��a��[��W���g��Y�	�'5P��&ފM�l�G耲j!����'�^��.�O io���ȅ�2"O� HC�
6}fN0�gEp�fUʦ"O��q�M	s����� ֙Q,F�q "O���nI3JE>�궠�0����"O(�0rbQYbVPY���^"�P�"O� 3d�, ���TnU"x��"Oz��p�H2��s�Uc�:�Y�"O�z�(�i�� C���Qz��"OR}h�A��mr
-�7(Њ @F���"O��kd��Y�e��`�8��"O�=���S��;S� �Op�|�U"OX�:%J�1y3����8pDr�9�"O��P��4<$p$�ޣ|-�d�g"Od�+2�ȉpX�}�E@�+$�"4"O �����*�Ĉ{?8M�"Ot��k�%S��BD�/@�0%�@"OѲ��ċ>�^�� �W1y^�0��"O��7 t�&�.��	��"O,`rJ���V���E=�"ؒ"O��20
�/{�4��bI�j��!Iq"O((b���
[�,Q���^ ��"O�����>	+ ŃEN�!6x�`�C"O� �d�@a��BGj@�֧�2_:<ks"O��"��Ů� sm\�V��s"Oy3ը\�tc�2��ƣi�d�'"OD��m�=�B�`�t(��"Ov��si�� ����A̿ :19"O`��#�Vzgf�3A��-@^����"O��w!ԝw��hH%�E���'"O�r�g��J�L����I����"Ol�	�"=-�`3"H�*$-���"O�x�7#[�� �c�Ai��g"O�=�
G75\�]c ��/&�d��"O��D�$�.ģ%��F����"OJS�0XM��FF �6(@s"O��X�$�?�zM
f��J9�"O����i����e+ȂP��q�"Od�y��V�ڄB`�X0NQ�e"O�}�& �
����7+�>(���,�y2!�W��S ��&-(��w�ک�yRº~H��'9�R��'���y������G�7"80�SΊ��!�<q�*�����'>p���E�"�!�$φX暭Xծ�%i�h:�M��}U!�$(V�|�O<O�hb+!�U�a����4��1P��8�� �+!�b�m�j�(��M��O��!�d�;p���`�q�($��ޕ�RB��'1������D�xr%���̈́ȓL���G�@6.ꐘaɉ5Md�]��uj�H`P@=2-����
�4@���ȓ/q~P���>���w.P�ua���ȓYT�Q�Ef�[�u`�� ��ȓawDD�l��j_=�Թ��r'�1Ga�"R��D�Vdh���"i�\(B�L�wB�E��e�c�<����Op"�X@�����:�DQ\�<�5�4
.ً�KLx�R�P\�<9��V5���%]�d��ɳWS�<p��,,�[DkW2r,�Q��K�<y%�5+��y�$�˦<�d��p�VJ�<Q�ܗ>2rT�N��G��;0�UC�<�0il_��;���� ���gz�<�$�Z9/-n�
���u,�e�@�o�<�`��0����0BW)uj���Wo�c�<y��˃l��R��:C�#PU�<�q�I�o~`j��
�y�]�h�w�<���Z�$���៪z��I�fX�<�D
6HH�e��#}�B}����Q�<�DC	%Ed�����%9ǜ����N�<��c�<$}��`�7�ʉR4l�K�<�7)=>�hؓ�D* 6���J�B�<i��B�?�ָJƎ~& ��)�x�<��c�� �*T��s[��"Bw�<�5O�a��S&^Ẕ��r�<��M��mP�	`��<��9x2f�o�<aEe�:1��N�	X�^��0"t�<�0*�8��5"·�3bi���Gq�<9��C��|1G��4s-r�<)#�/a3"�y�� I��&b�V�<���cI��B'��:K����MP�<���!:.�c�\.C��VD�}!��k���Q@�{�`=�GN̤E0!�� 6��M�6d�Xr��Xs�W=q!�$��4�b�94�N?Uqt�u��<[!�:wؽ��d���b@щ$A!�� ��A��uU��XE�`�G"O�`f�˧�� v��1Y��9FO���X�!:�Tq!��9�E����Vf!�$��4�f��q�lTAC�ݸ
!�S�6�b��4F�(Ʀ�1F�+d�!���V�l����+ ���3D��!!�dոkَ�[�oD75�VU�҈S�(!��_�.�uR`&vZX���-!�D��B'��{�f�;H�!�E 
a!�dK� ��Y�^= �A�݁~I!�$�?G�<l`�G�w'�D������F�DԅR�<����>v9e���y���*WHF�b4B��%ePSD��ybLۉVQ|Ly�jӦM޲�� �y�Y�(E���(Z`�&�yR`_.j�BDȄL�<"���R�_���'�ў��� Hѝ_8R5V��7�4�D"OJt�i�
a>I�� 2&2��k��V�'��}�E�ڐ"dː-G�jy{�K/�хȓgv�!G���B�X!ӔIMot�ov(<1�䅵t6��씱�N��u�{�<��oϻ��!aw+��o�!Q��s�<y��R'O�x(�"ᆒ8����GJ x�<��N�E�fy����m�1�lu�<9ĭЉ|ڄ��M�+�b�$��n��hO�f.��o�*^�e����9D�@�ȓZ��Y���#�J�(c(]�����(� �C�ze�dP7Q?US�m�ȓ2��ط̗
���Så�GM��ȓw�v%���)E��q�ר��g����O��=��%��@�&��(�,
��\F�<i ɔ�.�J��)��I8 ��~�<�T��vp��Q�&��h�`�s�}�<� A�"�d�uV�/|���&�]�<�SJ̻wr���6��wcX���eD�<��jt�P�a'�x����0%I�<Y,T�1�`.D91r�R��|8��Ez��"4��cG�ѡePp���y"O�aa$=�B��o�\�c���'�a{��]$g0 �b��;f�H������x��'~d����=uyrv�J�o���"�'�,���"P��V���cͤ��hO�H�+X�D���eH��@��Q�'�!����ul]�$��Q�B��	R��$|��'���Zw�Q>٠Ț�d�Z9�bn�'v@���=D��įۉ2D�;��M;r4�kׁܠ�M+V&�����Qڴ�~J?�̓��W�r�����B�;7|�� ��T�!�d��1�����Ҟ���Z7�j���æ��`��QI�yR@Ɖ>�&�h��\ �����6�>�J��j���*R��QcbT��4��4D�\'��6��@#1�Շd��x�ͱ�$G{��)�e{��*S�̔s�Υ�Q�
5p!�H�S#�@�!��+��[�CAV�IOx�L��cV6BN4�TaΦA�8H�Ć#D���nS���Y	���
�>M�!D�X�+�����CKUQ�,q�a>D�������ڍ��-�?hǴ8(��8D�p��n}�n���<-���aR�4D�����!��-�v���	�(y��3D�!�n�?E��"'̃��@�o<D��i��ӄ!���UZ�yb��8D�$c޵�xyB��­�&�BV�)D���6%A#DH�{�#F�:.�}X�#&D��(��s�܌��Y���i�B#D�� ���'JV��*uB� =�*��"O��H�GC�K���x����POHI�R"O�Թa��4k{xT����#*LE;�"O�AQ�<a��H1�,߃;�x��U"OX���JA\���KE�d���"O�(��J�:(�Ѵ�݇k�M��"Ot��2ʀ}w*QJ�*�#{/^��%"O����M9�<�:�����1"O��9҃O�|�����'�6,�6"O��(�H�RA<T�tf�
R�F���"O� �g&/@��A��M�n�x�r�"O����L�6��a��k_5iD��(G"OT�ZS+ݼ��Pī��z�\ܠC"O&�`
�eˆ���+�bYx�"O�]	MQo�����R09�ZL��"OXP�0��6hČ*U���"O)�І�-i��c����\�~l@�"O�E�t�\7��U�jI	6��%��"O��Sա�p���)EV좹�"O���_�w:�k��L�]���j3"O�`� ��>S[d�K�&��@��#"Oj9��*@ Y�E�1�7+A����"O ��LG�"zBP�R/E%�E2�"Ob�X�eb�X@I��Q�_�%	3"O�`���8h�ȼf(��,M�&"OB����
1�cB}� �{"O�%�kN<?�E�� �e0�"O���F����#%��|���h�"O�"D�J�`]!����dX*�"O\���#�A�2������i"O��y�(I84�,%d�7�	x�"O���JP�gaֵ�������`�!��(f<�(2�ǹ{h��!2��@�!�Ē78����E�ϔnI�]"��::�!����.D�C�Ԉ*T�W�C8�!�u��)���_�T�.x�TE�I�!��3K�$3uņ.O�&��0��*�!�dőm�`��ǅ/x��Ç4!�$B�"�thKW�9$gl�j���uV!��f�f�(�ŇV�Y��cT/S�!�D��)�Ј�f�U"a��Z���[r!��ۙa�b���ٱL�z���I|!�ӑ�r�P�ٝ�:�Jw䂠�!�D�#>�251"��v�:�[ʴ'�!�V4H�F����ҿ!�@��#]5`�!�$Z�!3�4H�ɦV�L����[�!�䏉f�%!�Q2ojP8d�N�!��׿O�Ba�f��f����go�[�!�D>r`M��Y�!�&@C㇁�
!�D938�xD��b�J���&ůd�!�:~?���ċ!3|�]��`���!�$Y`�@lC���Kn�%�D���!���})$�"K�&T�5�a@Ι�!��5ll��Ì�2Af`�Q��!!{!�ć���h3N@�[%�L��F`���'�$,���Ł�< *�(3:p��'W�( ޵L�I����9'PE��'�*8�e�r�D�x�J���)��'�Z�SՁZ#|��I� �K\�'I��`�(��p�z��$>NZ�B
�'���Y�AL�wl@3���mU��0
�'7��xs�ѳl� �ۖ��s�tt�ۓݸ'�F�Q"�)L�u��g�)s�& �' TL��l�4y� q��
>z�V	x��� %�Rߛn��yV-�3�ܽrP"OZ�S�,�.��׍.
@��T"O-z��3 �X��͇�����
O�7��8w�4��Q��HA��	�.'!򄄜v#�0ڀ�[
�|t���8 �!�${��d*sjS>��E��˩e��'�r. <OΔ F�C	(h*���"WҾ5���d<�S�S�x�=����(�4hň֢r�C�ɉSn�q,�?��[�'R4c�C�	�L�;SCL�l��1%����fB��j��Qk׍Gŀa9�胪k�,B��9n�H�+M�syh�r �`HB�'[ z��E�'s�<l{���?�B�I�<فs�ZP� <9�#]��C�ɍs!6q�E�E�.�
��cZ$Q´C�	x>�A��#�'C��	�u�?gɜ����I:(�Q�I��q.ޭ;�/W"J�nC�	�(��Tۖ�
}��m�dV=UjC�ɰ^���!�\�(L�@�`@��xq�C�I|\��&)*�x 0WAR�Pa$��0?�wFU���[ǥ�??��푱,Ax�0�'9x} �ɨOܖ���a��(��O����΁.n�Z��R<�g�Q5��}"���	���A��9*paR�	������7D�\��M��X�JUs��|YQl;��馩l`�ŞD��� ��5n������������<���Z+<�`��E�LԬ��)�G�'n�ygԛL�swL�8��������yA^&+8�i��Y8(��@�$��Py⍃�"\1�$ �0~���cƈwX��Oٸ���!)*��Ӣ���<�Zp"O�]Q�a
����-1�8��$̊��y��-JpiUd��+���Yd���0<)���ǌtS�Ȼ`�Z>��{��b�!�$��g�^AU�]9Y>��҅��u�!�L�/�L����Q(����B��!�$�L5Cw�R����P��3-pa}b�>� ��(��dW�C5L��y���V�<AO,Dl��Ru�]�40B,z��Zi�<��i��9��ty��'�)�Ӏ�P�<�r'��iD���͇,��J�&�L�<���ȗq������@�)��A@~�<a�F�-�֠�c-��n�Z�HRx�<9��x% �x��'�i� ��s�<q���$���g)�\��4ᄀ�q�<i�h],��c�_�/LD1�_n�<��7kf�sU���$a�c�C�<��T��ШI��K�f��Ƥ\T�d?�O�X�K�7�2,)7��R�^T�"O.US��#��d��/��x�tpj�"O^�X Ã�^���nM��f�c��'��OԈ���ӼWK�}��n�'�
�qQ"O
���h��~����7-_0M�*}���>�	�W�Es�&
>��)pjǪN t��	L}�N_����u�	!a�b�ٔm�&��B�	�B��UBEI�Wx�h�	�,+w���:�	>���$M�P�p@�6#�B䉞M/
88�n�l>,���_�.����$5��8x���)�Xr
u�U@�Eb�B�	�v����5L� dK���Biۑ\eXB�ɎsP�92��$D<��i�L�6o8B�	�_fI@,�39!�db�a�b��C�ɖ ��yq����-K0H5�_�C�ɾwphă�<"}�p�_/k�C�)� ~��uI��z`�Y���C��ɺ6"O�{5�Q=R�@�()M$E���W"O-FM֯h}��ӈ�5@8�!"O��cV*��&��D�j�ۀ	���'��	�\N�к%cC;�H)�����$H˓�0?ɗ�w��.������Qɓ\�<���"�2�K���XF|�q$�Z�<�$��I�R���,��L0�`�q�<�K˓Q��[��@O(ܰ�B)�s�<1p�\�.,�l�.R\f�
�]I�<��ѯE�D{W�ۅ:��X�7�BX�hDy�J�"�r�ۣ��p�H��`��HO��F�7 ᫶���Y������&�'�ўb?��C��G.ڱ��G^�X��X�6�Dh<�1�ʿ�p$���5~��ȱ�Jp����'�O@I���z�Q�0ۖ0
�Zd"O�ؚ$�I#@>��#�6��YG�d4�Ş~�z4y����,�bA�R�B�y,� �ȓL��9c�\3\dA��H�47�ʵ�?���1,OZ=���P���Cc��4h��)�'H�;%�Р(sE�/m��Mq���;-�*C�!Mv�#�dK)UbH�wz��B䉿q|��R)�+T4�B5��wb�">ы�ɀ5t�;�.A蝹�GA
z8!�T�#�"ɘ���y5���a��q%���U{�������$V�����Y	����F΍�y����2�ppm�&|~)0�޵����>�	ۓmi\�3��q�l�S�Z�z���M3Cɒ-5� a�a�Z>;�xxpi�'�a���N6?1����&��r�, 2g�ϝ�p=!�}�' Y`�p%�l�����Jߴ}�B�I�M���B���dt�aa@K&"����8��#)����E�S����+��E��j���>a0�J&��NJ�<��r��h򉎡HO�t䗔F,�$�<$�Hx�&�Ta��c&+ m!�$�:q��Y:wώ�,�P�q� #Z]���k�*��V�?����-F�M0$�$,�Zp��7�y���Y�d��Tc�=x����ґ�M[���s�p�R�	�$ ER�nۇ`z�ɣu"O.��ŅL|M����a��DR�"O�\ٲL�P���tH�N`-Q�"O�ab�tq��
7n�<� ,a&"Of}�%�	�"���Ql�_�LD�Ɲ�(��I�nC*;�бR�(�pfBZXFxC䉺~/�� p�-%�8Q�`؏Y�B�%\��E"ʣo�0����Cj`�B��x8�IbwȈ/lސR�k�"�TB�I�e�p�0$�8 +���$÷t��HO�"}��O�NtTش匷TS���tgu�<��ɗ�mX�	�(1� �)�VyR�O��Dx��1�h�ѫ\�	����	���y"d�:���H��<�@��ڳ���{Ӏ#<a��ą2N�Ă��O�W�6-��E�2a�~2P�̢*J�\�yQ�	��d��	,D�4���ڞ4]�y�G�h^�h* ??����$�O��"�3�d�Ol�[�"O�H�Ơ�<{��Ad�;WpXQ]�L����d�~�=���K�H�@�aϿ1$�s�h\)0�C��; ��j�5Y�ʐI�#G3����hO�>Y;�JG�q�(1(��$JĠ$|Oc���3��6O���ٵa�:N)�{GE,D��8��� *.H�5���G�<uɱ�4��nڬO�"���K/����g�FC�I�qM�D���§.��U{qI/ �$w�$+�Of�S�OF� ^�����:|Cu�J���m��"O
��b]�N�1��
Kp�r�P?y�'���I�'�(l���N�h���.E5W��
�'A����Z�����D�Ř�M���yr�Q�SMl���IPw=�1pq$���0<�P�I�n�E+D�ϛP5���Xp 'm$D�H�%�!%^r��� y��{D"D�4 C�Is�&�бL']���Q�d!D���Q�q��i�� <8K����"+D�4���ȩ*7j�y���6�)D���BA'xy�4�M=����� +D�L1Sd��p��S�k��V�d\�`�#D��ф�M,K�h��"�r	�-D�ȹbj����ƊJ�@"x(��,D�TJ���M�L$!"��c�8��+D�$���=���v�-��ɠ�<D����Wlk���e��U��-{e�4D��
m%c&<��7���}|�m;�2D�$��Í:��؅%�#�(���#D����Ė504D$�N�H���P�4D�<2�֒e_>��@����P�4E.D�d���,���P�-G�!��! +D��¥��4xJ��`�+ƞ@E\x�#D���f�G�Hl�@)A�4:x�,#D�HkǨF
F*KޤH'Ĺ!" �!@�!�D�W���䊣ld�i�N�=/�!�'K���W��1�tţd.�F�!��X8��2`H58AB��ϰb�!��Ê;�H�I=Oȡ;х]!�� ��`�	=<�ŉ�J�	n!��(�����d�ђөIG�!�d^�J��,��L��"B�C�7�!�s.N�¡��wx�	�1Rg!�D��%n���_�5sj09F��/!��T�$���Βe
гu��q�!�$A74����W�l�ބ���A�3�!�˗;9�A�ׇ05�<��tAӢZ���
<�q�f��Cr݊��6�m+�'`f��h{rl�ss�Q�W��ɋ�'~�xs,�gNֹ��"�D���'�=Z�.�q�|���fI;PX)�'ު���$�n��P��؅mD�\�
�'LP�Å%G�^(�Q�%p[&L��'�0���k�%!K��1��
��z�<y2L
:v	�
Q	����J6b�u�<��ϲ6�"ԥ��(ļ����u�<iuBQ@:����V5^`J���t�<�gH�<���oH(A^����Is�<!�@�0 �M�e�'m�����i�<�(�/;�h���VQ(�J���r�<��Đ�Sk��
��"����h�<Ɇ��&��_�PJ
�B"m�g�<96���9��,�V-��
�^�<q�)��|���śy�1r�K�Z�<�4)�w�^@�Y�uQ���c�<9A&Veڨ��ʕ�I�|���K�t�<I�mO�; PuE�+->���lT�<!�E�����HM�yO�)�ȊL�<����z��S�.��$а�KL�<��!D{���/�$��HP��e�<1@M�RA�QlѦ}L�P��I�<��Ĕ�T��AS��d!7l<\��5��}�$���������#�D;ct%�ȓ5Լ8�Ε�z&t��ٟ\�P���S�? t	 �môj䲬�W�<��}�R"O���Ь�.5.�9CAŉ4���c"O���̇�a�^�[@@Vw�\�0"O��RB�,Le����ݫ8���%"O@T1t���*,��m:M��� "O��� �̺w%Z��u�$<�Q31"O���l�(�"ybUD�&mv�!��"O,�V�A�;�]Y�P�$��!�2"O�5�GŢg�BP��*��0�����"OB�����)W��%��%0xz���"O��w�_�#��j2��<`�{�"O: @c�*rT��D���)��D�1"O e!5N�t�����	�6,�@�3"OBxS2*N��ɺ�H�'�n�Z�"O\�(v ��Ӑg��VG���T"OdC���%7�@x����I�B"On�9gGA�Z�0����ga�8��"O\���A~��e��\	c�XG"O�У�	�!�6bu�Y<?#���"O��Y�O@�c|<E�ҁ"Zը�'<)1R�M}�EƖB;�ȵI�!���w�ܯ�y�j�W��`ȕ�A�}�ڜQ0�I&��'f�Q�iܫpWQ?��HԊZ���2�B��m�Q.4D�������H�%CX�nR�A�p	9�n�ѯ)}R�JS���$��5��Ń?�"-J��[(r"!�P� qb`�Ь)I��a�dA�( �+r'�4
ǚ��t�'n2=�d$ʩ+�!
�D�~���D��qCD:):�I6'��x9���b�rIp��C��C�	-��y1w@Sb�z�Z������$�#�K
p�|��'�\��ë$rO2E���*e�&C䉩}��u�''G-�����ϔn���,݅ywv�'�d1F�,O<mI��ۙ57�}��B�p7�P�f"O���ᜀKYH�I��L�d8.�I%��:�!�4�Řv\a|����`NA 4�E��p=Y0�:k!��kqz�X '���\3"L=7,�1�%D��{c�R�1,�  �<i�`��Ǆ#��<Y��%�`��a�O�>�*�lB�OEx�*�&p(�'.(=Q��,�@}�aU�nM���RtX��dE��'ݨ��
�az�P��L�"�1��'�@[Չ�+s($E9�:UZuX�'�)������ �V�jM<�c�'�<�QE!��.,L�b�×b<���'�Fm�t �7:ΨH����#u���Z�4-�
�f�9�)���J��m��%+6ET��r��)D�(�7CV&-����Uz[BA(F���4x�-,o�^ԇ�	�bd^\[� ��v��Ȁk��Z34��Ɔ^�rȢ�!ٱ2/t���HҖ����T�|b^��"OL PnI�u���ba�#	Sl����	?=�P ]��Q>Y�SĊ�$��)�,E�'-�<U�&D���!PX(@�a+�,|u�p ��z��EB/��S��y������#�J��F�ô!���y����2��Q�a+��<$D���yR����ȉ�c�b����/Q#�
0�aH�b�G $�a|�*�?98�HU,�E�p�� ծ�6e+V��)5��j�N��P
��8l�݂��ɖ]�m��#�)�O~��iE;t���E%�/��1&>���덬8��� ��Õ}�v�>D����nѸ?[�i�lͼc�
l�$���^����eه9���m��O��#~�}��[�Ѵ8I%�$� ��ȓ=��b���*"���A¦Cȼ��S�~�����@6P��H5�����^�RO~̨�Ȝ	�^(��� Va}BG�  �.�c"�ȍ^&�;�J^�.�l�y�ĕ!dX�숥��0Q��~BH��0�X���*�RkRԘ1`�?�0<����P��b��&}��A9L8�KnI>:�
Q�"-�yrl�k~*e
�a<<�^��ņ)�٨��� <ܓ3n�9_f���9O� �$�#�Հ3����)V�	���"O@8�R��`�h*�ןE�|4�g�-"�,�Sp~�i���!.���� �����,fzșV�%_�a{��:��哴+��A�rM�"�~����F��Y�'߅)Ј�12�'�ƅC0-F�sv�D�RLE�xr��Y�}��d{Zw�A4W���CI˱��'=�"����P�Vl����7�6��ȓ܁r���L��t;�E�4P8�Ñ@+Q�&4�4ȷ2[p�IŃ|����J�q��U@�킴�´1��I�j�!��CK�X{7�U F�:V�B�x��Fȉn�8�Z�H�R��d{��eZ)���A�Q�� `�o:lOr)�*�F�Y��g���f��7�N���Ĉ�B�ȓkh5�c3���A�쓋NU���>�bS1rB�����]�8h���IڥF���T��63l~�rpʆ�a!�D� �"Es�:`G��"pɄ�E��a9R�ҥ2�
�#&$�/ �NP��>��h�\�Ո�DF\���br��`�<Qi�@^p�p���O�Bm�p�Z�f�PADE��|��'Ф��3����3�ٸq7�QHD�	�Y��̅�	"[M|��$ΏzWfG�g:LmW�� n�m���l~x�j�`����MV�AUB̫�A�-z E��D7\�eYA�b�S�}1���4E�O	>5`��	b{�B�I�H��1���x���宔��@ʓr��1��9Q�ҧ(��hzt���}����R�u��В"OT�3��fN�9���!U�&�R�Ep�dW@��}�D �����PY*���e��h��6K�� %�� !Q�(,��I�s�b�B� ��D�@<Oc�� �؋uV�PSF��64����s��$�����.��!֎�6 N��3'	��]l|��2�x�h��8q�� ҥfG-��1�^?�]�5Ҙ�#I����hh "C� ��C�I����g��K�H�T�@>%�q��`A	Z<��$O#6B�k�@=/�LxB&ʦ�˓2Uf���.�17��QЃ/*� ��I0GBv�+�@ˋ3��D��c�i@*`!5� ,��8[���-�b�FdW�!�ͳ޸�"��'��spH֮Z����b�x�{b���s�v$0���@�8�f���V}��x�K����5
�z���"삎_�x�%l�~�<YcJס���d�u�rY���>7�z=�����O�R�I�i״��;ê����'	���;��!�2�T�N��yS�߶1"�u��s�q֧Z�(K�m��VZ0�	��@3�~Mꕋ�� �JLI�Ep�����':4���	�1*�J����ό4L�
ϓ*�B��U�N�1Z0�2C¸k�6=��A�6*���CfB�SK����S�+�D�r�@=f�{b�X� ���h*;0ez%���*8:y*�E�JV��/Ѽ,�>��Ó'TU�D�p�O�<��"�&��9}|b<�'��a
ŋ�h�T�a#�b�������V�$��D�U5j�!�K�x��iM~*6j	�y�c̾i�4|��Qr�b���	\��x"ڢQ�^iӒ�N�X�0\�N���12E.�+���uoB7n�>�1i�#R�FY����06<Y�>,�P�΁	Z��y�c?8�dn �\��AB�@m:����L_�t� ��̻gu*d�OH�[a�'M�� ���8n̐*X�<y�,� }$�A�՛E����稍�%�~ȏ�d�J	^��B�-~B����-�yrX�W��M�����%��(%˧up�1*�&�Z-K"��R�hjO?�b���!��LM~J%N�%j�J�I֏FA�����#"�z|R�����~ �2иM��İ$��l��zQ)�.z���H�H����3� ̚ej�f�}���ߎJ��G|BF��]�X�C�,_������|a�U�5�>d��h�T�Ҳ��i3!�C��˟'�.XJ`�u؞�(`B[:r��a����6p�u8�jr���H�x�p+��Q�*��ۻp��m�O�7m��Nh+��ٜ\��E�l�.�KŨ�g�<ɒH��b�6��J��ZU�u��)� -�.� ���
��<ٵ��5:�r��B�a�2���\Z�i����"Nל��2	�A	�S��]b���s�nДS+���Y���EdV�g/b8��2Yd��ꈓZGlK�b�<1Ӆ�)X���5�6��2HZ8ˣ�(Y�䙃����#>IF	C	bs�T3e�<q�1A4c�`�0�( ���� xQ�	��C�.Xj6���yҮBP�X�i�Oe��x��E��f�ջw);��)Sls�(z&��<x�܄���'�<e�G���c���':��I���z] �Rtk�♛��#o�͘!n0D���[��b� �GG9"��h�)oӔl3��k�����>��ׇ��e<�Ͱ&��y�>�kJ8��T�'��+>�D"F�݌Sab ��q>:�s���.��z�3.8)�'E9Vk���ѫI�!�``�"�<��[G
�%��6U�uJN,h�2-�%%N�Ga}��ʝf�4��&*� 4kpO�F@X&�[WV~�bfc�HpT�T f�Aau�'�p��`�"dCІ)3�`t��􄃭uHZt��'�0�~R���b�c�B�:ԸT����((ȥbs!^t]�C��G�>I���_�<��$*�ɟ(cŐ��$
k�a��<I�Q�N�"�|�Ā�D��Ҕo�-x�")�.��yb��5��� �Y3&7䁘����dγgNj�	�rV�����H���3]:^i�ȓK��çf�)
$��%[BId1�ȓA�\��/��T/N�[�)��N� ��ȓN��8�"�"O^ӂOI'[�,��J��}{��p]��*�ǓOǜ��25phj��ZAR�AF��4g���ȓd(A(��J.,�dH��,�3/;Z5�ȓ9�
p�U,V!"��m��M��ȓZ. 労��.¬��KG�M)��ȓzpٚ2KR��&1�7��1v5�ȓy�h\ñ�KM.�T񓍖�!�@��XedSѯA�r�"�8�)�4*nH���sh5�f�L?`�L��[�3KB�ȓ�ZH0�c����Q@�4rR`�ȓ+6�M�@O�t�h�w�NC�꜄�R�.\+��Ħ}Ȣec�
F���ȓ#D����I@�K���)Gih��ȓ^�J�@@Ŕ�b��hD,�<3�v�ȓ�"��%�/~q���蝢=	�хȓ/��Q�E	'h��A��	~��H��G<�I��߿w��$Y6�	;úh�ȓk\<���ɉk-��Ï^����Z�	B�ª'h��(�"�R8؆�Q�U90!���I�w��h}^)�ȓ_s>����^�D!���Q�c����M�ܡ�c����HM��/YK�=����u
Q@g��Iq'�N/}�e�ȓ/_Z�y�O��jG4�)���	���ȓ/~L���)~��@�!o�(f,��JܚsJÐZ� �� �z D�ȓ`��Q�'
�(M:1��Vu�����m(�IiW���E�,)cŋ¿+�*��ȓ#�0�s��n�$�q��9��ͅ����@��l��c����x��}���95����d�3B��-��T�6\Y�L�k�����R�P��_���{��@��@�eE�u;�u����T��y\����K,*���ȓ/P�"�.��[�l"d��.y.\�ȓE(�LF-_�@��Di�Cd6@�ȓ{�la�i	+%1�`��M
�0"�ȓj�a�@��{��$�#.�ZY�ȓr��}���C�EtB<P�������dD%�'J�3n�R��?IDT�ȓ��hQ2jL�3�����]�#�x��m1��`
@�7��9@�Z&��لȓ;Ħ��K'yJ�`)�$ʓ���� ����p'�-m��]a�mF�{P ��e �x��
}3�(y�@�/=�R�ȓzr�$�BcĲ�ҕ�Wn��I��H�ȓ@�Ƞ� �������(��&s�	'�P�q��B�[ L���?9��i7I���<j���1�~��ȓ9��"!�o�B@���x6d��ȓ7N��ITVQ���s6��2�@��ȓz� x��ϼF�h�¥�E�d�x ��mm찢�]�}�XJ��V��u�ȓN&�5�Q&�NxᲇɅ�[5���S�? $x�ҩ��Ch�B�J� Uɦ�H$"O��HF�^� ��
h��]�d@�t"O�ۆ��&XiI;Ǉ�W8x%"�"O(1U�(Zϲh�P�2i?���y2JȂ!j����ĺBa��i����y¤�gL�! A( EO� �	��y)���I���$>���ð`I��yB����̍�\��q����1�y�J�-$��t9���Q4^�3��yĈC�l�� S8I�X�2#���y�T��d�q`n�=K�Υ��@=�y X,L�LAq�&��*��Ӈ�yb��d����HP�xDXP���V��y⁘�=II"B!�7|'�I���۩�y��U+b���؁}N  f/��y2ʞ.�t�
��%��$�L�ȓ�h�æR�DEZ�RTn>zIP��ȓ}Ki��M����L�w�N<�ȓ��y���$��=���,u=D�ȓ8��1��oB�y��9�� -{��%�ȓbҾȻ&aԯjN���# ��ȓ#t|X0�	^;~00q�C#�]�ȓL�@�d��/m������=���hR���R	i�<y3���~r�4���7R},�7W�H�$ώ�hlx)��O>i~�`Ɔ%D��ЂN�����Sǎ�C���Pҡ#�ɻ;>�`��KR�O���� �	� <JS�T;ے���'ln`�Ѝ��'ЮP��-����Ƨ
�R�rJ�;F�<�@.O��P��$[an(� ��^�<Q�Ϻ3���"�l
$�l1�.u|�{�(�)V�>���~�hq15ȝ�C�,Lp ôxH����P���^�yR�
	e:��f�/2�(�0+�9�y� ��m�phxVO),�@1�����'���#��_� /�eG�tdZGVX=Z1fۊ0�X� �dي�y�����d 6X8"�+Q�_hp���ώ���"t�Q>�(�>����*�R��U�� �ȓ�h�#GG�)����	��e޲uHA
=vNd<�B�P��.D�n�.PH��[���0�!\O4�vʁ�8�x�'�V	k��)����ӄB�B!H�'q�A�fW.}�����,9�d��}���Չ�ӊc� ��U�@L*<@ه 
'1,�C䉾��0]�+���`�h��዁����'��>�I${�JpS�$�V��͖{ufC�I%�Lh�($SK�Zm�RjC�QdQ`����E����5'�TZC�/)�z��>(�}�R�!84C�ɂ�6���(�<����� 7mZ&~�F0��{���i\�h�7h_VB��1�N��91����'_��k�گQ���R�
E�f>�s�'�z�*gN�#W)a{"�(�ܠ��W4���fJ%�0> �ܴ(W$a��`�d;���⩝�O���G�-_�8��Y��҇
#W�Ѐs�'x���Ex"�_4;&�$Z%�U�O
¤a���K�[�j )�	�'w4Q2����)CD��㤘�e�xV��$f�b	�B�j��s�4�w�M+T�r�R
<n�(؀�8D�<�#�҇s���!�$/�Ÿpx�t��^NTQ���'(�"���A�1p�.]��j��s�i%��P3Κ�bva�bA
�J��/�4��"���x�(ufY� �xG�Ӵ08�Ex2���'-\��1jL�!��U�Ѯ.�)�1\�@7��H�(�k��^#!��\<6��E[�\�z}�)�e� �v��K�H�5&��̓�_�\P��a�s�4yt-W�N~t���k^�dp�#�*D���N;Pz`8Z�G� k�W�LqY�7-���1H�1�^����hO�-��l��#I��A6a x�
'�'4��5:�� H}�eM�3s"+����S�0K�Ք]�j(��=�^��O3u���P ��h�(��I�z���S��G�:���.t9����`7~d�7`,CAfQ��mG�8�V�C� ���ӂ*�?pl��V��m'>�p�H?+�:`�S��x��y��)���!j��w�/h|xC��+v�@
���@��Pt�߅x�H�B7ˁ�2K��*��G��u�׎��Q��W�ŒPHr���Rǜ	H%�1lOR��#
X���4��z�*�k�Q|��B�3���NR9D�R����"������W���f@�#g�O�	 ��I�8�g�)�T�����. � ]�E�ƺ"��+�n���y�nŅ 
�A�٠���i��[&�Blh ����	�Pi��'��m��Y�da����X<��
��#��1h&D�Lz5��'Bbt�oA�!H���rӂ�Pĉ�H|�9��=�(p��i�\
� ��X��5��	I& 0��<Dxr`ߌGk�48g��^����`�C6�y.&�:u���N[V�&Q��'Cȥ	����X�|H���O�B�8c>���ė(!��]+��O'"�e*�!D�P�
��dE�b�� �|yQ��XX��D��,r�#@��%��#}�'���q ָn�옃!C�Y��\�
�'#R�at�=ML��⌓@��u�U�F�D���$�.,� 1�m�&�F}�ğ%$��i�+"M��`4���0>a����8��Q�ϓQ��B�˅�F���+Q#L��t"�e�/+�a"�W�\7�81�
��@�Ċ�2��Ov�`�`ų,N2��K|�tE�6h��Ԓ ϕ�M�N	Po�D�<i���"n�\����8pxܑ�A�zyR�
��u���G���6}�"|80��"���G.��dcPC�	T6�Y1DŢO�H�+�����PM�0x��V3x-'?���F�T7!}NIj��/\ta'5�Oza0�⋻1�r`c�
����,��P�NN�|��@�T�kЈMr؟���dʽt\�Њ�eǫ_�xt�To2�I�o��Ygǉ�z�$�e���V��Oo
X1�BE��;1$&�h��'M��a��h=zea�U�D�苃Q�Q9���W�)Z�JQ�ξ�H����3O@Ը$Ƀ526�HX��χ8(�B�ɔG�X吡����j�.G�w��6��: �Ұ� ��ݎ�Y���+���ɢHX�O��{⃄(	4�b��0
��<:�b�����~r�ǓJ]���E��/��P��o�>o!�DɱG���� ^�v��a�O	���SDi�I~h_�	^i���B̧@�]4q���p�ũ
�@�A��� LvPC�I%h(�����B�n�b]?S�L���<y6;T^��r@IZI����0��N�['�h��F�ZLz�ӻ�az���i'2�(�i�N?���Z�ά�g��Ԉ@���:!�V�p4��;��'5|��	q���� �@|�Ҏy�'��Ld�&AWyBD@�,�U�?���\1�"�����'�C�%D��ӫW�;���S�11^U����#?�nIp������mMCu~��|���Ǽ˅d�!O��M�g�DY�R�{�<AU���$�
���̚�^!V�R�U��8��:yΨ�'� )BQ�_b�'�1h�)T5bp������NM��0�F-�e�X�a�����R�僓[���pi�N�DZ�B�"$ ����"Ѧ�Q��\>h��oƬ��*F��]������>��ֆ)>�"�{3�v$ܐ�"O���)
>��sUʁ�*���3�	?.����>V�̀+�<��g�i&��0w��:�hɫ!���`܊���	0o��Tц��sT�1��/�M���*���F�+W��m��Ʉ��dwb�( %ߩk��:3�	�V">I�,N��5�:�S�Q�fd㲆�9��%(p�B;F˓24�p�� lO��!�V�6&2��ơɴ(1�9Oj�S���"5�b*�'	J� Wk[�db��'>1(qC��N�9��07��i�3�'�C�ɸ>�f9(dJ�h�Q����z��D�@���s��6�ĉ��I9=�h! Dj�=o��	���4�)Bp��;���@���r���Ba~�뗠V!ҳ�ء"�r�:G�8v������S
\��n��g}�Kh�>-�dX�?�*V�O���'�P Q+��҅9-w!4a�4��O�p"b�$ .|��Z�*�&F'.����S�*[z��嗅�P��k�|���X]jEp�'�z%0��O�?WB9�r�B�fA�)3�'j� ��T2)",�	�a�nPpƎ=U�� eK�S6J���)�l#4x�㠓�Q������ P�Ӏ�	7+r���"�,ه�it�c!�D�z<�kTB�"���X�'��kR������<9��56NK5H������/�Y���[��?a�-�k��U儃L��0⑲'���Ul�YS^�4�Q-C��{��Ӧ|��hx�y2뗇G��1e��Jȵ�7$�>ye�H;�r�°��!%�$�	Ӻz���~\�ɟ1��U� ��F�az�^"�6�B$�^�IOf�0g���HOz�ia�Q	Y�~)�'5���y�D���=x�H�R�ӱ%ǀ��RO!D���OC'H�ȥ��Ď�8vIJ0!�O6|�/^K��x�D���)2�'Ȳ��ѮL� �2\�G�U����'�U�q$�6G�a(U� =����O�|�pꒁ�p=��&�Tm��f�31 *ŋFE�Y�<����jp�0���ek��(�fh��d�x���VT 	�iƦK��x�ȓ-�@���ڲG:B9Eݏc�R�ȓ~U���LɄ1� ���,X(]��E~�]H$��,L� �4!߇"?\��m�p �aE�l�|=�cĞ�,�@���`�x�AF+��K��ŘF�Ȅ>���\��+#�ͮX����CI*n���ȓq�D���f�W�Ё�UA��V��І�UJ`��0D
7 �rCB� �&��ȓd�T��OR�"�y1!��,Y��хȓLDи�G0�%��#Ū�ʓ:�V=�C�]�BGK�F�W/6D�xa��Qs�����6p���%G7D������;�Xsw���(�A���7D�(;�"6^�*�ڧ䐻���A(2D�|���6D�,(�窑�
H�%J�3D������
+)�1�RdN}[��#�0D��1��R?,��D�
� ����%+2D��`2DD�`@)xw�j0���*O8x 3���-[�:�+I�<d@h��"O�ic�'5@\h�Jƽam �z"OR��G�X9+��H2�[U@���"O� �)U��<t���Q�
�`��y��D�slVБg�?��L�!��y"�@�c�
����,/��X�0��yO�&b�:�b�ՓŨ�����y���9�l��9=ĩ$�Ɠ�yR!� �*1&�0"�r��ЇW��yhؤ%�p�`���r��L7�y�#�9� �8��!	:�+ ��y"��<i�li�O
�2%�y!f���y��2*��gZ�g�R+��E��y��7 �I��P"Q�a�2/�5�Px�&ڃIښ��$&�-$����1	F	� ���C��\�f�Հ ������Ǝ{�ԇȓ6�~�b�O�8}~UClF �,	��a�XP�#O�	t|I�GgͦX�����^��9�I�<1���P�!�z܄�x/P�钫�.^l�J硛�~�(��ȓE� �� �6x4(0邆*�ȓ$��	�S�";
��)���p슄�ȓ{@&ՋC�P�f�i�+����Y���*�r7�9b����.ʄZo���'���Iz��?Yj7�:(h˓�9A�/���)�O�����ۃU���
K���O���j�/�.T��5��'��U��.V�P�JZ�p;P$6�h�#�=�Z�SU�i�,�����"�<˓T �9�`�^�|�toC&��>#1��8^i�YG 	
k)��x7ٱ�L��&u������wr���	�#B���µ*ʅ+,P��ޢ+��9*����\��X��"U�p�)������I��6�����I6Z�D���P�v��}b3���l�`o�(8���4��Q��� rbUr#�W �l"�KZ�i�jl,JoF��CM�t��iW}��rBP�j�Ɲ�����t�ا�
 &���I��i~.�S��Ov�@��76��u��-53�9�t��D��t�p��P�8�R#���Ok�3� �!�g?79�Pb��N6]v�:5�[�/q4�{��I�6.� i�E�*S�Omq�:@yЄ�/[<h��`<��j�CLJ���Ł)hd	���*&�a�c��_}�1�����*��0.��\1����'_l ��0a�R<����'Q���R���j�&�;�B��K:��,�/N��H:C*��ԡk�O����+07�5��j��L|���	�W9(�
c3o�TM�ԧL�@�Ts�����IRf}�,�Ձϕ5ʆL�1 �<�&�i�'��^�X�'����$Y�t���
��B��D�G	V|���Θ�y2 �:D�ĕ��+�=�PS��޺�y���T߬ �$EJ��BXX����'al%ӀcT0W�v��saG�Z�p)I�'���w�oE��T �v!(�K�8D�,��*X��qkc��[�5�+)D�ӷf\#L��86b�{��Ԩ�%T������$ܬ\	5I�	&�hB#"O� 2�
�m�L���T�r.�<�4"O�p�w�Sa�l�D/".�l2�"OX4E,�Rǖ���틶vo.в�"O�-Q��
�OS��b�kU�1l��A"O�V
��h?Z�b�J�DŔ Z"Od3FJ���qS��E7`�����"O����/�"H��Pv�(�(g"O����ZE�t Vb8&�F�$"O����̉7*=�B�ެ5Q*��S"O�6`	P<48!BC̒GbH�c�"Oޤ�qE��v�����?\8��"O�p��2����'�>&Q�lJ"O�I�G� ������žD�	j3"O�E8r�U�dH%�C�Dx pi�"O�E��KĆe"��b�@�-]Yl��"Or��"�0#�X��Z�WA�Ѳ�"O� ;����Hu��[�^3���"O�=�ӏF'WC�$ �BZ���U"O2��GJ0&��(��a8O趑�"O�,��Q TSz-XӠW� ���s"O��Buc��n���3i���ᒖ"O�i"��'ʈ��Pe�)R��rf"O�P(�]e�j��0�޷�v�+�"O���ӈ��xhx�W���Q t�3"O�U���R�3�Vu��MB=#,��"O��j� B�k 8�P*��l�r��u"O
AZ%͈�):�9��N�6���X�"O��ї�ԗ^]:A9�W�!#L�b�"O��$���J��x��W�HI�"O�l�e�p�B�g�ӓ� b�"Oh	
�$Щ���G��7V�0Q�"Oڭ1��ݹ1�,�+'lwFT*"Oh�T�_*J�,��d[�cW�=�6"O:��u�O�dՔ�f�АV�8B�"Of��	 �#s|�ԞdANu�"O��I e�ՙ6AR�TF"�"O��6H8�qC��4!�¡�"OJ<����B5\�A�S�p��X� "O�+�7\���B�J�wD�s�"O(0t��'ON�0����lY�qS�"O��k��]|�2	��(�kV,i�"Oh������!ԡG%����"O�$�c��:P�z���
t�"O���U��<>�TM����k�0y�f"O�Uq�N<;㎈(��.}b��"OԠQ7��>	��w��9obt�r"O����V$7�6A�$/L�eI��"O�H��d��}&N�"3K!8��I�"O&�ӷBCj*ډ�G,ܱa�>Փ�"O�� 7O��l�F��q�2�Y�"O� �q�/�@�\Ȫ���)D���3�"OT86 �:�Ly�HӋ~`E)�"O2��W��^�A#W	?j��"O�����3X	�e&ˤAk���"Oa���2�N��(��eU��0"O��X�c�"�hU�D�U�27��xD"Od��ɧ/���:cF��(Z�X"O���Ō�:{�̀�DG�P-�1BQ"OY����H�� ��eTn�E��"Oy"��4)j.��e@<b�^x�'K6�[5`�5U�"���:F��#�'��M�#b�+_�A�L<�JE��'�v��D�ȿ�v�2gfH�'�dX�	�'м�	Eƀ�P�Y:���({0E��'&z��bب}c��E�Т-��'"�@Cǋ<)���c�û-�1�
�',�	d@0H�q�	�,Oe(1Y
�'E��&�Ӱ!,>�!��$v���'jl��N��C�1{��V��s
�'����C�A���|����
�'��$���ʒnt<Kc���jY��'��T�����+SV�I��f&�y�,�#ø��ʛ=]���pv����y�$&]��;�@
_<
�i���y"*�.3[�ԋ@&�>U��0l
>�y�f�=f+�y�.���P /���y�K�5A�(9�g�ݠ�����y�Gϭ��0z3��'C̊�30�O��y�h��A��h�eς%" mJ�o���y�O�<�	3Vɇt�	�"���y���>֜�s%���xRJxs�Ь�yr,^-}��!��'[��\�j����y��ԥN��� �H+E��*�y2L�<]���'O�����IA�O�yb�ķX4���ӧNS
��g���y2!H+�>9�ˆ�J�rh�F�_��y�&�)a	��>��R���y� �NZ�Q�Ņ7�
 q�"��y�E�(r��8��I�!7����G��;�Py"�S�Q΂D�$ɖ8G:�Ӓ�O�<�G^�^&!bW*ѓ{��!S�Jp�<I��R�b�5S��[�M�8����	R�<�t��4#u���߭���  J�<C�ËZ6j!�vƜ��H����Y@�<�����:��}a*T��XP�F�~�<�Ą��`� њ�ռk�q�'�o�<�3I��0R��w#"T��0r��i�<1F☁IM<���g��ӴT���n�<��K�i|�h	' �PE�BMg�<9��U�x���X6�M%R$���M�<!GI�`Ů���1l*yz1��L�<� i�j<9�q#՟l� �! &G�<)����p|�0ME'/���x�$�E�<	c�ɪ\[~-���M�3����I}�<1��܄,L�eE'L��` Z���z�<����Ǻ���ן/Ӿ��C{�<���V\�s��T�:y����u�<y%)hKȴ1��۫�>q˄O�r�<y����,ߪ-q��	1X6�9�y��I	�&k��_݆�Ŋ �ybʄQ�P���a�*p�d��0�y�*ǔW�MH�*�"��,���yr�N3�q.Q�5}h͢����yB�������N��5 Ҭa����y
� ����bΘ ܬ q��C  s��X�"OH���.>�V����-9�Nh��"O��""/M�Y���r�ңv����"O\$2�銱|SV`0��O4*>4�C"O"���~�r �/��/���!"O L3c�|�	��;O �5C�"O����^�jS��I����� �"ON!��V=)T�*e�.��ل"OH���+Ĝ�x���K����"OU���a��Q��=��Uqe"O�%��B]� ���*�. @"O�`��摎+��AySn�+w���
"O����G�2��%nʡ{�h�ʶ"Ol%�EH�5~r�HR,Sq[���"OΘ�UEc-(G�ۭzDh\��"O���I�,(�f,z ,��h&X��"OVmHGLT-t*���@W�2��"O^L��X6hT��Qe���^B�;�"O�E�ߵlL�=��(ϣ�i�E"O.��$N1}zM�������"O�p��"\"�y�3��k�fH�"On A�U�3�b�F(k۾��b"O$��.BX�ˇm�/�8��"OP�Ԯo&�Z�-"O0}��c��gx�h� C�&߸�s�"Oɐ%�	�U9�A	!��w�f�;�"O�]�r�©a������Q���M�$"O �)�M�>؄Ѫ7�Ҙ-s��ڄ"Oh#ύ�S�l)�R?Q�4�"O~Mx���P�D%��G�_ff	��"O��GmI�v[`qc���-vV��#"O4�Pp�_�xTT�"��]kr8�J�"O�,k�� =�1H��,h��z�"O.9����"u�<�瀚X`0�"Ol8�!�� M�УBN�;BTl)�"O��I�`������s�z�`"ORA��/K7�넯� �P
�"O�2�E �JYDB� ������4"Op�B�i%ZX��O��N"O�sʐ�On��ud:�H�&"O~@3��ĳn�
�*
��ae"Of	��o��^��( �#Y(�@�c�"O�� h��@��I��'�Tm�%"O��CTp&q1�9Ȝp��"O��sv��u��7d�:dP�t"Od�Y�FF""c�O+i0Tx��"O���q��i�V阱c --fpC�"O�q��УG�@Y�0��S6��i "Oh�r��?�j ��S�8��x�P"OUa'IN�1+�R�Pڨ��"O����
� ���ЏF����"O�m�h5�P�z��Of�:4��"O@�YV+Ի�B����̸X��]@r"O��y� L�!�DiهA'��Y�"O
�D(|+�蝦H�������u�<7�U�V���PS��(�%�K�<7��%��011L�G�e(�H~�<Y�)Ϛa�TSfd��|��ѱ�P�<�a�ι;n���@\�3o~�!��K�<��'9�쩇m��LB�%�]�<�� �+�@�bw�i+�(vO�X�<����q�A�m�4"��Ѳ%ZK�<aBӬ,I�d"�LƖ:l���(�E�<�F S�_SHM�0K
�RX�9��D�<� F�L��W�1 ��FS����"O��P`���(�R9a@+	�K���`"Ofy���G�Ft��`I��J��"O��(���g�0���N_�i�Ҭ�"OB��L
�d����OD���8�"O$�R�d�xZs�?E��E*�"OPբD���2*R�00�ǀ��,"A"O�W�R ,Ԥ�"�K�8O}`�5"O��*3G�uA����Lӎ"�L� `"O24�$��3z�� ���j���"O&P۳�KY��!/�_T敨֭�O�,V��Mcϓ�M����ު�dB�9�v)jVV~����@�=O'f(� /ݻSP�ё�m�':�0if��;~�3
�TB���hR�^����P�`��G����]� �$x�Qb4��'�0�8�e��mzx8`2M����ݴ����͟PN<���?�L<y M�l��#� �_ P��n�@?���t��Zdむ ��9�ߧn/��K�z�h�O�m�?�'����i��7�W60�	A8o21��H�;��x��'�:y���׿2�"(+�����L̃�4!D7�AD�0�R�$��iE~r�W�`.$�+&�S,�1zG�
�`&��b�EL&.�rt�q�8EH�@���-6��ˡ�+�ɍ1���D�O6M<T�h��F�>QJ���2��M���	wy��'}�O�OO�-�D[3���"�ɚD�� �'�����e�6��m��e�? �bݩ�N@¦y��Yy§8j6M�O�c?)�A� �h��`�+mTL�A�x2�'V^|���%���@bR�H����C Q�4c�&���Ҧ{��=� ���'��8� ĀX<@��s �v�,��.�h��A��ϊ�]A��/tBb�4����O8�d+��~�]�I=�Pے��i-�!ru
� j�'4r�����1b� aB�R�d4�[��P����d��]�IL}�cN+t��4���Wh��aE�f9,���KJѦ���|yʟ�b��*� �+����*
�~�is���4 ���±�J=�H���Ǔ+ct��>��ӫ��d�
۴�R	׃+?T�qQ.��:�4��i�7�����eI�'�4�*�c�=�fD3S��Tdj�1�C�6���g���Y P`#�?���\r剁������Oǥ�:A���a��Xw~5�F䃯\��$*�� ,O��8�	 ���I��WѤ1"�����ʟ�;�4���O>6-#.�҈�uFל������
"n�����l�x�4n�rB ]K�ǗSmP@MX�N沉a��S�Jp�A�gT�7�n�����r�#>!�@�B5���sg� 5����.�5cL:�B˔=t~x���r�����0���1EB�ig1O&�p�G=6r8{��/^�0P3�jR��z��	ٟh�ݴ�?I)O���.�e�ԄܐF�Dݸ��C��qOj��D�J����NJ�iЦ�y��
W�$!��4��c����O���<1�lP��4�M㛢r��L +D+w}��K��a8���	,9�E ��:�$T���P�>sN,���!E�@-w��9Y࡙ a�8]⑟ ����&Y-N)��@%�h��f�'�J�i�.``�9s¾|Zm�Q��N��%�?�����|�	�x���Q��d֜�+%(ٝ6��0��^ܟx�'o���BY�p��|�T�h	׊�:;I�e�3� &��݆�L5�r��[��j(�QA�lW��nZѦ��I���ݴ�?9��?�L>��@9�P  ��   �  P  �  �  *  :5  o@  L  �W  �b  ]l  zu  .|  r�  \�  ��  ��  v�  ��  ��  L�  ��  !�  ��  ��  6�  ��  ��  ,�  m�  ��  ;�  1 { � | �  w( 2 �9 v@ �F �L �M  �L#�靱I�8��tE*���"O�$��L�'bj�����΂<4��ش"O�Ȩ6���U8�	���& .�1�f"Ob)��E�z���q-�"O�(��B�\n���ФV_��"OL�!��� ���Ja�I<�[�"O��R.\?`����lW�=zh��"O�}@gL�`��R�B�
0�]Y�"O����o�-vY��'�!["����"O���Kl;z,
�G��!"@"O*|�I�E:d}Ar���/���F"Ov����L#0���ҥ;����"O�M�R��D��\��8�l�J7"O����A�Z�z���N��A"O�D��-e�F��VA�3���:�"O��`IO^x*(b�� .h<24"OP!��l�CVl�#��#L@@�"O�m1'bȅl�� �P#��eU�] `"O�Z0����s�"R~9�r"O�@c�e�"]���1Q���a�ʥ@$"O�i����b�h5,Rz4���@"Ol8{֤D�����rdO���r1*O�!cA%%��[q���n��	�'?H �gA	27]Tj��M�z�6D�	�'���혶T�>쩷E�phֽ9	�'0��N�{K�u�#��cɐ���'��(���8����d�cܳ�' ����_�?���B�
���
�'�.�S�/�q��jSd��9��A�'��S#Y?	�T���܈�*�`�'��T���;V����X�5�Ji��'�J�j��F:���&^0����'�8��$	��P)j�,�iʦu9�'�"ř�.�<[&C��g�XH��'R��"ŋܭ9h�X�H�R��I��'%���e��h����V��3�'�Za��a�v=	@o�8xuB�'(�}k7�[62�����/2=��;�'Z����� �~^�j����{�PE#�''N����6��Aևs�0)��'h��7��X��"'�4n ��'�F铰�#E `�XA��H�JH	�'�Z�CA��
]q�@�%�_O�v���'�hx��L���q�:�����'vR=��k�"�S�F�/?ꀁ�'�f퓱��<=�p0���:�&UB�'\ ��Øb: �eNGb��'{�`�Ȍ�O0�*�*�W��H�
�'���H��	�KS�� �,Vf� q
�'���v�\ |A~����͐S��,R�'D|(� �x�x���"S�#�m2�'|ܣ�"]�Li"s,��ʜ@
�'�nAaV���#$�h`����c�'��h����Z\�a�ѣ:¡��'�;�H"@�� _"�0%��'ޘq��ھX�� R8�B��'��(��ĩY���Q�)U|��x�'U�����¤0a��+!C�a8���'wd
󪈪V'TU����;\:R���'�����.0��j��?(�̼��'�² �6~�Ȃ���#�! �' �r�._����)�.Y;�'��T�4�R?:0��HC�,w��s�'L�t�ņ�쵌�a�xYqר��y
� ����X�'$c�$ʼ#~����"O*%0���.f�\h�"ܫdx���"O��IB
L��I�����&��0"OR0��ŀRBe����t	�#"O�Cp.��In�9k���l�T��"O�	��΁,�ބ���E0CGtqp"ORY��(��%搡D/9RP��"Oj�д�³Q����F=ILn��G"Ojq��-:�2�¦�0N��0�"Oz�Q�29�P�H��X� �{3"O:��g�?{��x�W���0�"O��������o�❙ "O��'�R�uk���i�+9tv���"O��'n�JdL ���Nj�[�"O���U@�+�\�#��@PjDTd"O���π&���Y2��[���K�"OȰ"C+ea�\q1��BaO�A�!�DU���ӣk�16�ZD�r@!��ڭ7]�&�U�)����+9 �!�ĕ1��̉+]�:ZI��}�#�'F44 ��� q��r��K-{�P�(�'xH�Y�e�#Cı���̧�����'zN�2���4kl�P�Jٖ �dq�	�'czdǕ��\�$�I:
X��'0�(�Š��n� ��\y��l
�'����2EA#<{��s�h��'���+r�߯�z�쌽}u���'�6UZe�x�ܚ�C�)�ͨf*D�x8�`D�;K&8�f�NT��) �*=D�0	�n-ڤ�7�K7��.D�$��U6%�4b�b�*��*�,D������&l*u���A$LhH�.7D���@����`� ��s�FD(�;D�\ɒcL7�ܬ0@��E���u�+D�<d�:a��`'�J�2Ĵ`��(D������k��z�b�Y�Ph�*%D��������Y��H�lZ^��!(4���W���n	���^�a�� �BV�<���H �H��U���Y�|��f�N�<�V�E5��I�E�ҷD���iDc�<t&p�ƘYK�-U��b!��^�<�$�!yR,&��sg �K%	A�<��@�jP�Ձ�X4g�v�S/�v�<�ӂ
�2}����/
p�;�I�J�<�R���l�q�U�t���X@�<i���`�xs�R�Ty4����'b?���AWKvaY��R�u��Ց�=D��;���	Xv��$��@)�S1�7D�����޷DM�1�S+�-��]���;D����	Z�0fn[<3\�X6�>D����m�B
�})q�c)۔�E� �Q��F{*�@���� $�6���H�w�xtʥ"O��K�ͼ[�Qd�X�`y3�i�Dx��s� lY�j��G] �!a	�>��"O��cR�@�5:��@�B� ��t�O���$�DpnQ;N��=y�Ɩ�B�!�du�j���.V�Q�0�p��o1!�� �kH��vc�^�ބ�3'��b�!�d�����`�B�2Y��f (�!�ؕ��0��(��b�X
�N�E���8D{����8S������6��f����"O� Z��k�����˗-<�0x	7"O�E��/m����4��.Q�ҩC�"O��t#�\�D �ɑ |�����"O� �|끅O�`$N�񎃓R��Q�d+�S�'\��u�d��u3<�[&�ӣC��X�ȓ \� ��1^X�J"k:��'ў"|�D�ki�!�7d��	Ѹ�"��V|�<I��]� j6��V,��xV8�M
^�<�wO�?P2�L�A\�J����2��T�<)%�
DĐ]K6�H�䀊��W�<I2�ŲO��{�k�)t� ��F�w��0Dx�K��+���蝔���ٲu�<��K�.:�f���^\tP�Q� v�'��y�C�6*�| �We�/$���mR��xr��tr��׫��aHd	H�!�Ē*6�1p�_6D[6�1B؃k��y�	���8�OΚ^j�eB!1|��p?�P�M�Zz���GO�E�Ȁ�4u~R>O�O|`����O+��'���-�2�8T"L,:uFA�'o�����I�� ې����۱�y��iq�@�f��V�%�S�<�O4�m;�	k!�J�ˑ N�$4��'���AA�Ƞ�c�Q�$p3N<y޴;�D%��M4O�����0@� ���1=��h��'���-e1���w�A"v[��¤��0ܜC�ɝ�P 2���9&�vЊBc�0W��hO> u&�%d��xvh�9W�A�6!+D��q��0%,�!N�X��}Iw%;��:�O$!h�W7 �P�#�O%6Uʬ�u"On��Ѫ�,x���N'bh$�T"O0���Q�&�*���+E}��k�"O1GCE%<�j)q1*�iؚ��"OT�8��ܙ�R\QgN(Gd*S�"OĨc�O��B�P��唽HL~���"O�|�qᛠ!��|S�d	$"1* t"O���C�%]��YCS�0�3�"O���S��t���t��/����"O�̀Dn|ZixBͮN]\u��"O�Y���
&Y]$@���0"����"Odͳ�1%�����OX95���s�"O���oÚ,��`��N��W����"O��Y�St"`)zu��
��S"O�)��F�f����V:>� �4"O�H*�F�4_��`"JG�R�����"O)��ʎ�4U,���n�s|,�v"O����B*��}���y�q"O�tg�BWZ��1)�x\��Za"OD`�`��$���& nr`s�"O��gR�rn�*`d
+h��"O�<I���9* J��r�ǂm����"O�b��`ZXq�p�[pd�B�"O��:����;d����� [�U��"O����MU('�.-���^=RRL���"O(��E��P v�8��^Q��a"OT��o�X��@,Q�7\(; "O��r	^
�p�f�!~�	(�"OP���dh��c��X�D�"O����� !B�.�:bO\�x��t"OF�ib�(UN(�#E)�]+�"O գEhs_�q͆0S�x��"Od�2�'��1PdQ[���%v�
�"O�i� J � ��-h�bL@�"Oܤ��ui��'�ޣ�q�v"O�E�Ηpg6�	j�t"O�;ÍH�p����Cχ�6�rt"O�嫓�;[0Ut�7��t�a"OЀ�$�5#�^��g�T�2�"O�=��ɇa�P� ǅ84���!�"O� (�C��Ù.Yʕ���	(��z�"OL�2F`�1��ء��%<>2�3�"OD�b��K�6T9�G��R59�r"O�3�lNצh1�/S�>V�%"O�prZ�7�r�yPj��U�)C��'���'��'m��'���'���'�@�鵄Z�N�(YV���~�(e0�'<2�'�"�'���'X��'���'�Ii�e:bk��#P/ԇmS
��'1��'��'��'02�'�'k�m��	?��(�zh�s��'���'���'�2�'�B�'R��'�+�P�F�ʱ��)#Q�:��'�2�'�'���'���'K��'��c�,���	��!�x�NMH��'��'R�'���'���'�"�'�,��F��b2루_�7�����'�b�'���'��'>��'q��'Ӟ�P�+.b'j)�\�d8��W�'���'�"�'dR�'O�'3��'�t�9�)��bK�iж3��QI�'d�'`��''�'J��'���'j�X�� �;���e����4���'�'F��'b�'���'�2�'��R�n����W䍙Lz��pf�'cR�'~��'!b�'�2�'p��'m��3
� K�����X�6g�@˥�'�B�'�"�'���'���'m�'��� �n}�ի%��J1�MKw�'��'�B�'���'�Ҥk�����Oތk�!�ƭ���Ƞ+�����Ɉxy��'��)�3?I��if��&��T���S�\�p�DZ����S�e�?��<�(��}��'Z��(�mҞj1����?q%X��M��Ot�Ӧ��L?�`�U��B��v�$K�:�Ɵ�'��>E��U8K��!�+��|���צ�M�u'�A���OIZ6=� �vj�3kt�� ��Dnb|���O6��e�Xԧ�O8�p��il���R����K�l�H������Do����i_b�=�'�?�j�+�0�UCc�}�����<�(O�O�dl���(b��gm�\V��nC�X8�J�~�l���ş��	�<��Oz0�Dbc� ��Ѡ��Vl�a��p�I�)����f�$�S$)�r�ϟX��i��*tAH]&��IB1��EyQ�L�)��<q�l׆d�|�ba�Q�>�����k�<��it.u#�O�yo�`��|��$ѐ[P�5 �76N�bw���<9���?���8B,	ߴ���n>�`�'DC1�5�+}]�c8A|"�{�0��<�'�?9���?���?!��0���.'
E@"h���� )O,Tl t����ɟ��IW��ɟ�;�A�Vx���ݚ(a��0$/�)��$�OV�'���J	%�F�i��W�x��B�Rc�] !�w��ї'�����I?�M>Q/O�5�U���K�0!��Zq��R���O���O��D�O�	�<���ib�PC�'�Hh�m��
�Z����� o`�Qɑ�'��7m=�������O@�d�O�t��"нvjxшu��a�F0R�O�'87M1?�H�0\��}�S��5�W�ցD��Af�\��qAW�~��Iӟp�I؟���Οd��S*�.�d�p��ղ3���2"n߼�?���?1��i>z@�'W�`Bش�����3E�#��Y����q�5!H>����?�'j8��4�����=�S�C�eB��ʔ�]*(����X1�?&D9���<�'�?����?!�NڼYy��F��G@�A�s�[��?1�����Gɦ=��O^�<����ЕOB\}��
��s x������4n$d"�O���'"�'�ɧ�)��[׎A8��G<��-�2gΏB�@�tm;Q4DT�����S�v��'�z�	�fBmI��Ӈ�Z�D���G!���	П��I���)�ny",a���QB'>"����!�Z;`���晁0�$ʓyc����\}��'A�!8%�ٙIr�@ǒm�'�r��?0T�f���{vc�n��~
q�Tr���Ui�$[��Xֆ��</On���Ok�i�b�'�rX>�9�\��\X�1��!���#e���M�Fދ�?9��?QK~2��7e��wrLݢ�e�4��0�`"x>�%�'�|��D��Y�5O"��������l�P��a!9O`z � ��~r�|rP��ҟ�AU�Ҥc(�ڃ(�19�8��P֟(�	��x�Ihy���"�°Y�T���r���H��Ԥ~@i"�#g�8%�D�	����O&�d:��^�7]bUK�J�g�bd�Cm����>N�=�3��A�M~��砟��I�^����	��@�vI+�5������	� �I]��y��1wX�(Vg#-��hd��0pSb�jӪ0�%�Oz���I$��s�� 	�t�&h%C
l9YȠw�x��柈���$P)mn~2[�C0x��~p�m9"5-��lҧ���=�M>*Oj�D�O���O���O���� Bp��Q���RW ���<�`�i�l<�bP�t�	W��LAP"�=w���X�����tXZe���d�O���2�󉔸x� �;1��D�)I�R�#"���Ec���'��lA��?qN>)(O���b+(�fС�#� '@E���O.��OH�d�O�I�<qg�i"���'=:�)T�bl�᧌&b6���'7�0������Ol��Ol�1���vlZ�cԻj�h��nU�9�7=?��{��'��!�K~��{�? �6xx�9�b�vm�9Æ=O2�$�O��D�O����OP�?A8e���.y.P���� �oYşH�	����Ҕ��ğs�4��|/l��ECXv�Al�?Ҵ%�O>����?ͧ1�ݴ��$�;�2��g�%:���)ư7t0<���?�~B�|�X�T������C�^��2�B֥�_s������	fy�~ӄ��o�O:�D�OX˧bZ� �0�O��^�"w�ŝz�m�'Y:듲?)����S�TNZ9��Z�@�
�.����\䤕 �7F(���<�'���Iz�I�d�(���۰}_��xc�J�6PT���ɟ���ß��)�Ey2dӶ�����~�,�͓���Tꗔ]z˓a%�F���M}��'o��
�d3(B�3qf��0��I���'A&K+ ��� �%��	�q�Tă��y%���� A%,i˄1O���?9��?���?����I�B��(�M�-"D����+�Pql�4ض��'�B�iZ���J����/�c��,��o�
=�IΟ�%�b>Q"t��Ѧ�͓f�@���	�m����CA�!>�n�͓Q{�P��I���%�P�����'���P7�0;\8����@�����' R�'\r\���ڴ>C�����?���B8�Q��`��ɑ Zx	9�bJ�>Q���?�H>���'_���� �#}�e"���v~r�A�G�:��g�3��O�8��	1B� ��d��L��wX ��&�i�Z�M���?���h���$��Sh$�;D��#j�z_ zrd�d���ȵI��ɛ�MÎ�w�vQe�s`$��FťQ?�'�Z��I�&��)�'`T�U��?QE�̛'cj�pS�Jː��ąI���'��	�����ڟ@��П���A��}���H��3!Q�l�z��'UD7m�˓�?�H~������d�5AA��E
 �p�T���V��I̟�'�b>�j��[�R� d�H�5X��*�aQH,m���V�/����'��'E��.QXMG��L�� ��w*���ş��	���i>]�'J�7ML�|���p��LH%�<"�r���L�����	'�����$�O��D�O|p"AaÀEn��ȧoˠ!�"M*j��k07�1?�4�(�@��M���ɺAe��o��͘�H���(s�\���������	џ��Ja*
�I��ِ�Q�{��H��a�-�?����?���i)����R�4�ݴ���m3�)1F-��B�"ˡ/㊍�I>A���?�'}�T0��4�����r��	�eA����q�W�Y�tϖ=�2H� �?���8�$�<�|�	���cW�F"6ZQ���3%t�Ex�h�d�;G/�<������	`�����j�
�����k��������O�D&��?�Q�[�(J�E�
HadJȐ�ՌQQ�AFæ�+O�Ȫ�~��|r悌JJ�T"�j�,�$p��9z��'�r�'���TY��(ٴm�2̉�I)8��m���a�ڵ�Ǌ�����)�?��Z���	�Zmjj)h��(F�Ҁ��矘� *�ӦE�'��[�`J�?	��D�څiĉ���A� ��,�p�V4O@��?Y���?Y��?�,O���$-b8J��٫]±���O�ʄn�tC�$�������J���������E ؑ59zYҕCG�NSFq˒�Ģ�?Y���Ş�T�޴�y�N�(����*X9NyFt�fO��y�
������������O���Y�.B���e\/l{��A쑲4����O����Ov�m�6�S#=���'��B^0�N��ߣ.e*T���ѣ|.�Ou�'#�'a�'��$(&ŋ'��|��jS��� 2�Oy���'Q}ڭQd��Χ�?dD�O0E��!x7�HP��;� =�g��O����Ob���O�}���2�����? B`!�ȝKH����G=�v�Ή,�r�'i�7m1�iޕж�9b��e�0`�6hK�d���I�,�	�L;dTmK~����P$�'{b�$@3|9>���Ä@T��O>�.O1�1O6�"�L;&��t���(�H
ƚ�<x۴wZ��(O��D(§?�lr��(V���˞�'�$�O����O��O1�P��c�x==��"L�Ljj��З7�.7�syB�P�m���������䗦U2�ssCD�U L��7���-����O�D�OR�4���\P��of��nӰц� �5{X�����)�y�z�*�p�O��D�O���L�2((�"Ei�6[�|(ӑ�R�:�X��&d���J�^��M�\QJ~"��&h�y���.�����N_�^����?���?����?q����O�H�d�:@�IP!W=R��PEX���ɗ�M�#���|��Qߛ��|R����ƈ:�R�5��(���ڪE�'������EB9gK����P`�"F�)��4	Wk�tj1@g
?�����O~�O���?����?��Q�^���S��3ƅ�!r5���?�,O�Llڑ0@U��䟨�	@��JY�bT��=}�*,1�O�9�!�'���?I���S�deʝO��81��_� ��
��/rW��t��&${�m
�O�i��?��1�DR B�rq��H�o�$�1��G�Ӹ���O�D�O���<�6�i�0E�E-G����EZ
a��t۵Iޮp\"�'�7m7�4��H�'��@��l�: �H�	fL�(!R�'� ySB�i!�	5��c�ԟ�S�? ������"*��:b�J�RY蜀V4O�˓�?1���?����?)����	�&;̔b&%c�,!d�]�h��n�-B�ƈ�'�B�I�˦�7w���֋#x	�R�c�B��	���$�b>`#N�ͦ�7JZ���1�=1�M]b$�1Γ.����O�%(N>)O�i�O��@�����D%V� s��O��d�O>���<�%�i�|r��'~"�'�ZȹL�	;�%Ba(P�K5�5� �|��'r�듀?a�����1�S��5y���@��P�'�DB�a�+q0�:3��� �ߟ�:��'��P�qhS�wLj)�5NY�L�J���'�"�'��'��>�0JĪl�2d�AƠȲ�+�e��8�I�M��]��?	��B���|��y��]�W ؠ���3%i�,�riמ�y��'	��':����iO��5���ן:�JbjU�7Ā�4�H�4E��r��*�D�<����?)��?a���?A'⋛/c�D����VNd($k�:��D����J� �៼��ԟ�'?牱i^.`�c�8�l�F@�+��@�O��$�O
�O1��!�T�0�Pq�O�h��%R̀7�r ����Kb���o
�`Mj�IByb�M�ZFL�P�	
Uf���th�l��'5��'��OI��ʇ$�̟��W�L$r�r����e����ڟ8��4���|JBP��������ɳ`\�h������P�A��3%#�!x���Q�'Δ��V�O~r�;dl8� \>z�����A�\`���?��?Y���?�����O_���g.@�J��1`s*�#%\�����'��'�F6�͐9���O�ioZ{�	�)���cE�2j���Ƌ1 ��9%��������$�o�e~Zw�p�� ԯ/H�pRd�M�0)Vc�B�"
"�Hu�	byB�'���'���4f���� GZ�C����$�^��'\�	��MS�"_��?����?�)��]�ҧϔA"� � Y�+��S���i�OT�d�O��O�Ӥn�CC��Q�2�
w�R���H��" �4��mZ���4�L���'��'fa�b�sV��p��*L�1r�'1r�'�B���O��	��Mc��#W�q�Mן:0�5���Oz�f�(*OP�l�l�?0�	埘S�(T8m�����	�JQH�qP�៤��9U��lq~�N��5|0p�}
4h�-F����'M ?z匔����<I,O���O����OL�D�O�'^B�bCdP#E,�A�DbnJ���Ȧ�*c�by�'��emz���G��@� ��H�U�L�+�����O�)擅P��HmZJ?�o�!�`�#φ�|�����|��k�N�;��X�	sy�O+��8|n��K" �Ѐ`���v���'���'��	��M�[ �?����?A��U�w�4�cbO9f
l�w/�0��'��듗?������h�
&-��d3�@�D�2)�'XrȦoӳ˲MR���N��dR��'��)8�дP"0��Đ�	0����'4r�'
R�'��>����7���� ��ȼ1��� 9�������M���7�?9�8|���4�d!ɅA��
Ų��;M�iZ�3O��D�<)g͟��M��O��k%&�ⅡՅo�)	��B�}�q�M"Z0ȓO�˓�?Q��?9��?������bkBiUҩi`� �P1j!�*O0�mZ%SZ���	֟H�	u�֟ �t�O>{�0��W@)-��ea�����OH�d<�󉘁.ԡW��(�(gи?�����tExʓ@�JT�c��O��K>�+O�nA.��'�݄=gȋr,\����O����O��4�Z�>���g�x��!���2fC�+S�	�d�k�hs�x�hC�O���<Y�EJ�#��M)�.�"�����
�/V���ش��$�*K�Bd���xS���P�3AڐE�;��j� �j��$9�OJ0R�Õ/r �4)�NS��BӲ
�<���k˛`���צA'�L��� ��	�\	R��cGݡM��'2B����܌D�F��H���@Y��w犔y+��uC�^HHI���O6�O"���'��pe��`����eȻ�2s������e��dy2�'��S� ���r�۟�Ɣ�0��8r�����؟���n�)�"̯&����Ɠn���ClU���+�'a�7�Uey�O\<���M���� ATl�bWZ�a����?���?9�Ş�����3����y��QaR!(o$�WG�#���	ٟxڴ��'����?��f�%���	�c��|�$(�@eƊ�?I�$yD�!�4����<���0(�*O�Q���<R�>`{2��W��0O:��?���?9��?1�����:�́�{G���3�	:{޸m��zB�'C��t�'�7=��ru�i�L��C36Q�P��Oz��$��ǧ-6�7�h�X	C��6Rj4t����Mt�}3",r�l#�B�KE��2�$�<����?��MƁZ�p�PK�_���1*�
�?1��?i�����QP�gO��8�I�2GM����)�tc�j��!�qcHh��ǟ<#�O��D�O:�OB�#��L8�����g�!(�~l ĝ�`�UB�-W�����GZ��(VB�ȟ�Ѧ.R>I�lD{��W�|=�$ρȟ��I�,�����E��wF8�YT �7e�LI@��%WoΥ���'C�6S�@���O<n�S�	۟�]*uI���p�՟=-��D��)Q��	�����Ο��(Q����u��(V�4�*� ��ƪ
u/�u�DN�s���%�$�<y��?Y��?q��?)�Ƀ6O���8ECO� �xk��� �����A��ʟ���䟔�Ru��R�m����zXI�&"9~d��ԟ���u�)�;%���.�<	���STF*z�z1��b�ۦe�-OR�S�k�7�~"�|�Q�<�bL$�P�
�EƝ.t��a�`������㟌��џ�qy��m��+�M�O��Q�)+��{�|�����?Q\�(���>Y��?���u�`�
�Ŀ(檁@�k)T��0��_2�M��OR=����&�������wPz� g&�y�%[�BG�HҘT��'g��'��'{��'���]��c15g�,X$	� !��{�G�O����Of�mZ���'06M6����iFIKQ���`W�a�B]�6*�O��O��;w�7�6?�d�\ e)��r �`*,��Oݴg^ ��Od�	N>).O���O����O�h��GBGu��$ᔁg��e�O���<�U�i�����'���'���c��X���;J���#W�Z���\��I埀��W�)�*P�t��a4I�\9�Å#l�^�8`�Օ�M��O�)��~2�|�&�ym�"ᓨG�l��E�?'��'Y"�'z��T_��Xߴ~kl��b�Y�Z�v����4@��t�"��?���-���$�O}�'��yJV.�~=����..�dMk&�'�id �ƛ��~)����,.��Ai��Y���#F�j�[BoȃU�<�Xy2�'TR�'9�'�R>������F�{*�}���0VqIm�1�Dܗ'#�	O���ݪVk(�j @ۇS#�E��.
�-��ğt$�b>i�K���̓+���ҡ��[)Ш���䰜Γ�ա�
�?�.�d�<���?y�#޸bs�8�t)�p��A!bGM��?���?�����ZЦ��7�oy��'����1�SF|�\�P�R�Q̭@#�|��'�등?����
}�и@#J� ��!�������E~D�%�pQ�`�i�������'�M#5�J�����H�TE{@!3m2�'�'XR�s�]�蘌����ĳon0p��B�Ɵ��شB�V�P���?��ixɧ��wN����D�>XC�&ÄO��*�'(��'o����h6����0�/?��I�'�j���DB@Ĳ����30�F�O���?)��?i��?����k� :���je�4~�Bhh/O|�nZ�d����I�����]����(F�N�%���j"k6.�9Id���$�OH��(���	=�p�wɝ6i��<w��ggP\�P�}w�I%b�Έ���'��'���'O��y�'��-�v)��%3<�%���'Ub�'R���T�@�޴.�8Xi�.��a�c
ʒ��o�'Y��[.��\O}2�'."�'�p���.��9K���͊"^n���*�	6��6��p����\��D����<Q�3�G��@!a$�]5h���:O~���O��$�O��D�O��?A���P�C���BGE�u�^`���Dy��'�7V"��S��M{O>�t(Q!a�,�K'�F�F� �(�����?��|ڔ�� �M��O<�U�}���i�	Pඔ�"c�'N�����s��O ��|���?q��Qy����&NzɂVO@0FD���?Q,O��o��>��	�l��c�4�p<�ղq��FIꩈ�e���$Na}��'��O�S�d�<�:�ͿT��4�'X-n��HV�ð/z�J�IPAy�Oʺp�	&AL�'Ƣ��!l�+�H��0bIoܨj��'���'}����O?�	��M�rH4>P`��Ϫ^W��J����� h+O�m�S��XW�Iҟ�.���`��Ԩq{>7�Z�?��z���Z޴��$D�hHj���O��ɍ6�W]6-Eha�Έ?B!�)�'H�	����il�Ɵ����x�O���xa�.�Ġ�Ј�8Z ,觬y�l�:���O���O�����Ħ�7m`��y�L2j$�gKeW
��I�L%�b>�@��榕�TLf���l(r1��N�����!�^�y���O�8YK>a.O��$�OȘ���)ZIrI��_F'�,+��O����O��d�<�U�'9��[��?a����".1*��-Z�枫"��`�2a�>���?II>�t�S�s���g*ۈ�# Ot~r�T��><A�i1���tyX�'��ar��+O�W�t�ǆJ�2�'��';�����:����g~�yx�!	熙I7�A����4���,O�QnO�Ӽ3^Y�-�p+�.o����÷r&���O����OH��g�s��ӺS�dA7�*n��|��(��C"g�� ����*3��O�ʓ�?���?A���?a�>/$�s���( 8�+���)�*O6HlZ: [�H��֟�IV�S֟�(զ
;�.ђ��ܭnu|�h�����On��'��)� hQ2���I@�X�~a��m�H��S�-(~�ʓt��5�D �O��H>�,O���GGȽ!�t�:�̅�Et�ۗk�O����O����O�ɡ<AA�iބ�µ�'�R����.�)fMV0����'E
7M$�D�OX�'b�'���XQ�F�@3�O�ڔX$o��Y���i�i��	�%tfe!&�O*�l$?9�ݑ�i�Q��*TΪ�2�ھg���f��x�p@�74�a�J��bAU�P�"l�'�B�m��-3�?��޴��Ob���7
ħ#�}boN%(�p�L>a��?ͧor�P�ٴ��ē�� ~`��4k��q���o�P)�EE�~2�|�R����埸�Iޟh���U���k��U#
�Z`��H�����py"�eӨ�*B�O���O�˧e�����C�9qج�f�I���!͓�?�!V�D��ڟT&��'Ku&�RġW�f�洉����b{PѠT'��``��(O���4������9�`�O2͂��{��Xqլ��c���ڑ��O��d�O����O1�^˓i���H���5m&4r�1� �1qN4Ya�'��Fu���ȭO���VP���)7h�UH|B�i��#�l���O�!�t���/d��b���D�O��iY3,��Hʪ�!��A&Zp:%ʝ'����������<������IZ�T��.>v-�5	Ũl|,p��Q�n6�ź0�,���O���<���O-mz���,EǠH�`.b�5vOMߟ��	T�)�S�VX��o��<�uG�aאQ0�iS),F��;1K��<v�>��[�Dy��'�n͙V9\xcTBÅKA�'I�)m���'r�'��I�M�����?����?�2�R<{����ݬ!k��3ǃ���'�^��?	��N�-;J�%cǭ�Q.����^���[�"����W�=rJ�������r��d�0
!J�c�B��p:�
������OB��O�*�'�?�P���"��!6&�@�x`���?a��i�xi�$X�1ش���y׎*�������n��w��.�yb�'�R�'�P�(�i��	�[�!���O�D �1OT�n�	�i�~�1���Wp��~y�O9�'���'�b��d�A�TL�!|�����̷_��#�M{a�>�?!���?IN~Γ+J^�7M�;��ABP���t��W_V}b�'���|�����5��i¤��s��٣%_�X���U�ixd˓-��"$䥟�'� �'2~آ�@� �Ћ3	�!V�fm �'���'�����Y���ٴDm���Y*pIS�ؐZ��bdK�=0����֛F��Mq}��'���'�][�#ԼcN���_�kz�	硌�QX���L��$���������6	��L�2�}��ͤ�?O��$�O���Oh��O��?�@�َJÎ���k^�ż	�kV̟����H;ش����'�?��i��'IΜ5H��Rc�qR�"�U�\ �y��'"�I$Фl�B~��L�P\�Q1D/�U9��B7v.�|Ja��T���Iʰ�ă�"=�9`�)vr�8$"	 XuT� �M�ݠ�`�x���䇇�!�<����<~�� ���1q
��ALκ��2C�H����g-��[�q�'�������fϘ�Sb*�K��ЃHX�]ʃnѨu���P�F�;\�*�(Ąޢ2�.���.�C@lmc�)��\p��Ze��?1�41�K��Rkq)��c��-��BmŬ����K� �Ꙙ���%s�pM�<��t��,��w���B6��e�6m�U�.2�٣+Y�R�0��o֛eS��cF�Ē0��I	Ц��Iӟ��I�?	bF%et@��7�Q 
����îZ	���?y�$Y.`Gxbҟ�����-"���vI�<�B�Q�iU�IaE�P��4�?����?i�'��i�):�u�h�$��`���Ħw� ���O�E��0�IRܧ]j���D�4/΀��錔P��n�?r�*ɚ�4�?���?y�'=���Yy�$8f�����s3(�ӵ���6�-L^�X����|~D:T�@�:*�1xÖ�
�&��i��'nR�+y������O��I�m �	�u���*,��']g�b�˷�;���d��ȟ���ʐ~�4�䤁2Y�8��&��M��9��0�wV��'��|Zc�F`����+6��q)��}8����O�X�U/��O����O��4��1�U̵�L�(�iA�d��xaZ�<V�	Xy��'Z�'���'��#r���@�X��D�5Q�(A�V�'(��'v�X��Z$g���d/<k�:���K�c�j��D��M�/O��$ ���O���FL�����J��<�7n�H�(��%��|N(��?���?y*O���)�|Z��TO��g	�-�F�/)�nm)�ib"�|B�'cn����>�Va�$wL,�F�^!7����l������؟ܗ'���0l�~����?���0��{W�^s�V�"�L�~{"P �x�'�R��t��O��'FJ���%[�=p2L�FY�7m�<�&
Ɠc�F�'O��'����>���f�xs���L��KdKn�\m�쟔�	�W����?���4O,�R<�� i�Ht����M���8ӛ��'���'���	:�4�`	%-�9!ip���$I< &�ź�/Ѧ��	ş��Iy�)Γ�?�sNT=D��8`B!H�8��QU%;���'�"�'�Xɣ�'�4�Z�d����P!07C���۫%�`(
�$e�p�D(�dLJ��'��'EB!�q�91g	�)�`��gc�$B�B6-�OF��"e�l�i>��	X�f����D�hhjC� ��	H<������?�,O��D�=4:��'�@�qfH<
!ã�<���?Q���'K�DI�Z����5A@
6�|����D~Λ��K��D�O^���Or�$����<�쵓7���!Ap��kL�(�p]���	ҟP'�ؔ����'��]���/t:|01j;R:t �f�#���O��?ц����Ou�e��-?�����ѝ2��t�O���U�?����D"MK�'�Vt����
y�^}"	�u
rmjߴ�?�(O��d�j*8˧�?�����1r!
q�_���Y��E>W���%����Ky��7�O�ط7����E8
���W$�e[��V���I��M��U?a���?�*�O� �2%A�$���C-�#,P��iZ��ܟ���1�ħ���%ie�����?(�b]	��sӌ)�0c�O��D�O����D�S�t�ϰn\��F�.%]\��C	´t��O-��Fx����'x�(#ԉ�.FB�8�Tn����DsӴ���O��ŸY�Re&��ڟ��JڶD�7��'^
��˗-A7u�Tnܟ�$�0�����O����O�D �F�%T����a��>���
��
ɦ���� �K<�'�?N>rIǲ!� Q��H�_�����2�''��|"�'m�Iٟ�
P9�萪�-
T�����3���'J�'��O��ķ�����y���V*���	+]W�&�3��'�X���ɨ0Z���T�$u{�.�+�P��A@�H�*pm����B��?Y(Oԍ�Ұia�l�R�Z�\��uaPQ@�R�O���O��$�<� ���Z�O_��C1A�wH��#�ïun�kAsӤ�D�O���?�*���d�|�"�\j�h�s!��X�2X� G������'x�Iş�[�@u���'���5�Sq:��G#�$�)J��L1�ē�?Y,Ojeq$�i��K�O�u�d� �z��h���c��˓)����i0<��?	��dO��>F/���T�Ke;��5a�.��7ͥ<����?aǞ����ܴh@��H���(jV~���a^��=o�����4�?���?��+�����ŚG��l �(̓rX���&D(SUb7�OB�d�OܒO�s���I=0�R��c�X
A6�ZǍ�,� �ݴ�?���?a�
�n��&�'���'���uw�Z7��5aI	 ��@�i[��M����d�"��?u�	��L�	7�ހ�QA:f�ࢆ\����޴�?�)�~_��by�'�����؆;>��4IY�8��ܫ�ߖPR6-�O�Y8!7O����O��O���<4������r�\s&]��:}'hԫ�[���'�b^���I�h��1�l	SH�53�����
�k RI�3p�x�'��'���'�2c T��6m��C���B���~�RS�A�a.	o蟸��ןx����|�'_�B1����($8�x�OyW�	J��7-�O�d�O��ļ<9���_������� ��q�C�k����@oӂ���<����?�o�µ���4eF�z���;,���cǐd�mğ|��EyR熲�H맏?�����qj�~kp\�d�	�o�Np[PD_!N�I�x��|�a�i�|&��'p(>؁E�:B�h5��)
5:�n�GyR#R�L��7m�O,�$�O��iu}ZwX��2�f����ur���b{0@�ܴ�?��M6�����ϸO�00��l�R��AJ�	&U�@�HߴF����w�i��'=R�OH���F4Y�y(U�8.���A�Lpuo�+[�4��4�'���䚇$�l͂���0'����<A��m⟸��П �����Ĵ<	���~d� ���#$�7�zpS�#�MJ>)rc��<�ObB�'�"-g{¤�PA@ ���ЈQj��6M�O�y	pa�Y}�[���	Hy���5��;HSD���˴n4���B������A%�D�Ox���O���|�*�2=3�ᅷK�Y���X��L��#�3?��byr�'m���������N����� ��<cɘ��w�����	ʟ�������	��'[T](�he>Q�2���h1҈ꥫ�����p�˓�?/O��O���Ea��D�,	}s�l��l̘�@ӯK�{�|m��8���$�	]y�DB�f$x�'�?�1 &I�+�":M����ߋq$�n����'�2�'�//�y�_>7MUPa��!r���5a]ƛ�'gR^�,Ҥ������Ov�d�`H��lһ(&����+0��a�PNc}B�'�r�'��邟'��^���������-�\����٩f;�!nZYy򂟜$H7m�O����O��I�i}Zw�����+6���_Z��۴�?i�q�.8��?�-OD�>Q	��ҏ[0���f�3mȀ\�j�6 ����Ʀ��	�����?���O��Q����r��Qu��sB�ɸu;DhF�i���?I/O��?����s�6���<j6�,+� ��4��4�?���?! ����|yR�'&�Ą?s�u�G��}"�1Y�k�+כ�'����)���?Q��sd ��':,�^�0&G��M�#���?D��q�	sy�'-�I���6H�4J gI"��0���\B7M�Oސ8E7O(�$�O����O����<ys%C�H����15��sV��5�2pɶT���'
�\�����,��~Uʵ���UT��Q"��x�uH�Ir���'5��'�R�`B�^=���cړ2�d�C7�H�J^�xq�U�����O��$$���O��$-��$I��ڝZ��(T��X��͆�0��$�'���'gBW�0(��ޥ�ħu��)��`�w�%~��U���i�r�|2�'�bOE�8���>�J��58N�n�$\R���ڦ�����L�'���r�K&���O��	H�M���P�d�)-����w�\�ACM%���I��K`l{�(%� ��j���G����؁b%�Q�hmZxy�,Θ+v�6�V�d�'��,?yb����y�g�(*i���٦9�I���J�E#�ڸO�U��A2ph U�6)���Z�4\Ӱ��i��'��Onc�D���C�#�������H�V%���C�M��j.�?M>��D�'I�t�@��	�S�ύ)���s�n����O���L7e�R��>9��~
� "Yu,�+��!q�gV:R��|2��$���D�<Y���?��Oj�D)�努2`r �2��9;���ش�?#f
\_�'P2�'�ɧ5�.��0X�L����,���X��Ky���:�y2S����ϟ`&?yIgkN[��b�ϛ�)�8�!��Ա��}��'��'��'^t zփ�:c�h| �ib<���FB*_?�[����ן|�IoyB�(�"�S�X<*�J�%C� P&K�B�OD�.��OF�$őQ=��D��3�Z�2�`�}*@���l͕#I���'-�'!�V�L��j���'V�t�"�̑�f����#@+��ر�i��|��'��T�m�qOdI�q�'n �܂倘�y(���ix��'��D�&x#J|���2q�/e���dN�)p@8��)X��'Rb�'/��v�'��'��	ܨ?A�,��g#>j�0aŽY5��W�pEO�0�MWS?����?��Olj���8x��� iD��i���'���`�'zɧ�OPZ\)um�X7���2�E�)�t)�شXu2��$�i;�'��O}bO�	L)i��@���.�f�"�l�@L�'b��i�Oh@TK�+[f�eX:����������	Ο��ʹ|���I�O�I�ؐY�ԀQ�1�*��FLG�,h�s���Rh����x�I�dC�O��:��$�?4q:%�p&���MC��8'
d0��x��'b�|Zcd�2�LF
)�x0*p�R�n�l������O��$�OH�A�Ȕ����6<�Ց�/�
�ta�@��'��'�'��'�N�{&��<#��s0`i�QC���'3b�'��	�� ����͟LkW%7FH����a@A�DdR�����M���?A���䓻?I+O�YPe�i�pq0��#�ڀR��;��x�O"���O4��<!��$i�O}�$)��ƴ�#J�3��T�Ec����:�D�O�>1�)T�c]f�`�
�Q!�AWæ���ܟX�'n����<��O��)V� l�y�B�(L��0 ��_��d'����A���c�ȝ�Vd~l��41��YcuFc�˓/z@�i'4�'�?9��w��ɮ9��) EՃ,��y�J�vպ7�O����A>W�)Fb�U�ʍ	r,�Nv��"��yN6��O���O��)I�I� ���	n�l���]�BLZ�Q �C��M�gOI[�'{����(�����;�Hd`�%T�h�P�oZ���	ȟ�����ē�?���~�b H���� @�h�ܲ%�Q��'��u"�y��'�B�' �����B��X�n�|�z��Voy�R��� * `�'��	ş�'�Zc�����aJ��y�g__���b�O�H֐�������I˟��'�2��Z��[W�J+K�xAIvf�cѮ�����O�˓�?����?	�j���b��>l��8*���^m��̓�?���?����?q)Oz����|"7�@-�)��_~��RaN�٦=�'Y�W�8���`�Irt�ɂ���#�!^	����YZl�r�O����O����<YUg�+u�����f�w���s�ڴ���� /�M����d�Oz���O��8:O��'���bD+I�F��� X�z���X�4�?9����ץ�.��Oi��'e���z�����"��
���£���b듕?Y���?	P�]�<y)��$�?!�N������Ush�Ѱ�u��˓'���v�i!2�'�r�O)h�Ӻs!�L6B����c判gEX0u����՟����o����YyB�i�7AtRtX 
	1:�اՐQ��6 E
�B7��O��D�O��	�h}�_��#埅�X��V.-6�)iT朡�M�V��<�M>�����'Y"h�ԉ&��Űg�ȅjWN��s�����O����M�0l�'���,�}����4�O�Jf�]93CW"�lߟ�'Ya(���I�O(���O���	�2_=�8���K%��VH�Ϧe��)I���O��?�*O���.� �H������c *
	��P���u�D������	����	Dy�K��.��V�
�]1B]sh©#�`����<Y�����OX�D�O~�C�c�g�|�	���vd�"�rG���O^���O��Į<ͧ$��O4�Y�c�U�m�A)Q�<J�Tqݴ�?!���?O>)���d̗e���D��H��a 16$*�� ����O���O�u(v`���$遟,vRp;RaR�e�B��/�k�6��O
�O���"�et��G��Z����$�>IxYm�ݟ��Iay
�2�B�J�$��T� ��^�����:{1R�4�\Y�����	�0vF#<)�O��u�w�u˼�ē�Ti�4��$S��HlZ����O��iRD~2��%��Q����4���p�Lʏ�MK���?qLL�'pq�h���$�<^���Xd�d�(�%�Q��c���A�<�b!ME0�D�Уm�Lq��?�d�A6��aaǀF���� ��!�$�(p=x�G�ЫX���{�oO��5��նt�0�*���AծTk0�_<d(��ƊեDׄq�lH��ĕ���<EZ��5�o����ր�,٤�a%,Q$1Po�#q;�m���N(m
���sݎ!rW��8��!���O��P����:m��`���MLv@at�Hk*�D�O��d�O�P�;�?����`ܴ�@t��cqu��o�/���I�o[V��o�(�q�0�e!(�U�ӃS��%*3x�j\�MG_K�pa�'`����)�)�t�����6s�O�!�� fq�`G(KK(�V�Y�%.�	Jb�O�&ړ��'YD�T'K����o,��	�'�^�K��ײt����S���qC�yrl�>!/OR�����x}��'�X�B�oD�AF�J��Z�dl6�'�mK�D�B�'��i��&�h�Hu+V8Y�������Տƶ\̎M�RF�[��e��I�-���J5O�8�]S�'(D�{��Mn��Â�Pd*�Y	�5����ǟX�'%>rc�ʙau"��w�Q'C���y�'��(f(Q�mR���A7�\X�'+
7�pȕ�æ�v$ 7��HyZ���?O
�l^`�`�[���	G�����J��mZr��ciD.��(R�4t���'��hAQ�0���Em�YT��T>іO8���J+	�,a�c"D�"tzI��g�
#s�
��u��t�uF���H7?6�t���ʲ��c����ɒ#����O0�}J�nn> �%̨A��lhF$�J��ń�GXPZVґk꬀	BE��%�ʅ��	�HO\��u��2�9g�܈S(&�:t�h}��'�⮄���2r�'R�'��w{�!���V�n�<�C��?C����V�
-��e��.�O@����xz1��'�Le0�=y3~����A0Ke��	s	XD�`���O��� Ǆ�����d�:c�'0�L��T���1rt=�����D�9cC�ODў����؜���ĩA���cC. D�0Ӣ�ˤz��f�@�Sϒ��*>?9��)*)O��� H�:�2l��(��g����#N�K�`�`�k�O���O���˺���?��Of��5m-&a����J�╲�ǃF(<�����$PLH��o��(�)žj�B��	(�=���3Pp�![�6��B���O �$;���O,�?��y� bH�5@�!��}4`B䉴g��|�����ġ+�k���Bb�\ШO��r7�ū��i-��'�$Q�Bfψ$0� ��G̠��@�'t��jt�'���tR�|Bm�=[;,2�-�a���U����p<BN�n��2���Q��.`M"ů�JnV4��4���d4�ǒ^�~�rboG�gr��g'+�!�d�h�� �烨p��H��W.8�!����A0#	�=k�ES�L��kJf�P��/扣�ƽXڴ�?�����A}4�ċ�}Kv|0�>�� ���6���d�O���G�O�b��g~��&�����Z�UѪ�R��Ǽ��$y�j#<�rV��#z�R5��� *8��)�-�R��٘AP�����&1�>��@�U&��
*(���+
�'g�B䦟�xL�@K�	�Q�[	ÓH��$KDmU6e*x[�"�u�&���	2�M[���?	��"c��I5��*�?���?��Ӽs�ȏ�k��p��K� r:�΃$�z��%�Bh�4�iS%�b���y���xRKL�9�=�����:�У7��Eӄ���%*>�^dc��J%�	(����xR)q5L�w��6l���`��^1t6��O*��X���4�D�$�O����O����=�h4�$�$�$ɢ"iƘ+��C�	U	H�ZC�;G�"ع`���zb0�	q�����OxʓA	 �����:~]\��IH21�"�ʣصnIܬ���?����?�������Ol�S�W�d	I���J%4�3A�\	Rؒt���:�02���#V��sbÉ|
A��'�2C�I�!,ɫ���:ehta0f�XCH�O������f68���(!�Ty(`͜nu!�d0 ��D���L�|BE��bd1O���>2�U�ay���'�G�!4�\�Y��֜WM�b���RA2�'WZ)z�'�2��u d�xӀ�O
��T� S2��F/ޫ+�t}x�'/Z����Ԛ]^"a��_'���6�����x��Z��?�����dxi(qñh�%�d�B�Z}���O8�4�)�'q�ʸȗ C�z�
 K���-8����6���¡"۬L�`)W�n�)b�,�y2^���D��5�M���?9.���QB	�O�T�&A�r�䠊qJ��*��a��O��D�;/��d.�|�'a���
��������(~YM��Pq'�S�'1*�����eNH��gM.��m�O����'V1O�� Q�n��x��E��?`�Q�t"O�U��IK�(�,�T�)Wb���'�L"=Q$�Q���]�#��P*A�#GD��'O"�'�n��  ݝ2��'����yG�M�tu@��oX:""��˹U�u+���	j]���-�5�#ɜr ���bBYX�8���;P}t����؂eX�:Q����'ΰ��S����I�� Ԩ2τ�CrX��d�./
���G/4�p�w~X��#LH>a�E+�??���)J/O6�s���0~�T)JΦG�d�8���<0�z�#���O����O|����k��?9�O���#�#�<��-:F����Z'�xR��;�`Q14f�+o���ꇬF	W
����'�hQ��A��&A�OB��]���ʺ�?I	��n�d�� �}�XXc��D?&hN�ȓQ��l�U,�!��<��.�>�`��<Y��;6�A�'�����5ضq�E?f�|D��fV�r��'��`��'y"1�͠�Bv��ġ��[�	_Z�Q�B�2����l�8s�oԨ�p<��N)9��R�I�g϶͉s�^$~$�\�z�4�"�J߭7 ~��ēD?Y����d(���@c�|�L4�ţ��;�1OB��d@�x0�r�^|��a��Q��!���Ѧ=�q� Rc,�&IQ|:U��Av��'��ԡGIr����OzʧZ���*�qn�H,�l���9�,U!j�R1C���?A��@��?��y*���4h@$�%l^F��H�r(��L�N�'��Ű���	ǀH���&MY�s&��7�H"*�1�\��R�S��&���Hr	�+[��0+�h��%�х�r�d=Xr��/y���b��L=X�@<��	-�HOFA(!o�Y۶�߭4Qp�*����I������)���z�-ݟ�����i�q�����;B�ĳYB���5��.�&��#���=�t&?c��bL�;иl	�L9b�
0L
LV��"i�<A�ċ�=���>�OzaRl sMh̊��PUf� �&�O�XlZ͟�C�Jџ�>˓�?1�f�{��kj�k��h����$1�OL��3��#iL:�W��-(i�>�ܴ��f�T>y�'�&�i L�	b�$��@	�N8�ddӻ�x�0�'�b�'Vlqݡ������'n����R�E�&���D�C,QX+�(u�C��mArLQ��U���@`I!`:ŉu�+�Pq�k��=�t�4 &V�	�:?���'�O�#HJ�*�,���[��=��"O0;P�BR4�MK�c!8�,�W��^�Lة��i�'�i���C#����K�I?f���'�J]�	�"�'��iR�{�b�|�b_~򉺧m�xT�{4FK�p<�5��o�j���"c�G�e�w�W#�@ń�I�0@�$�Od�F���9D�&kO+��	ot@�ϓ�?��������Q�� %���0�݊9=��ibO>�lZ lI���d�K&�6�ć2'�	Vy�6M�OP��|�!���?�4���8��� �P)|� �[ *V=�?��
=�%������0���3��I��j\>�u�� }���3�O�`���	�-���F�SH�.B�>�g��H�<�"\ u�t����|�|�H�v�<aBƀ@Kn�+��B'P���PMY�����dˏq�N��g���~h��1�l� i��l�h�Ißp�c���������	�� ��P��6����d��	�n��<��l�Cx�dв�Rfd}�F��	=#�}I` &�I&�v��d�=hL$��h��/Lr(+�]�l��c�4j�Oq��'��|�`�6A8��L]�lҽI�'�v���	'�ر�H� 9����OLDz��I]-Wk\�v�^$�uK�A�j:�;���������O����OX�;�?������
͐lz�Ia��	�k\���/��w�~��'=.��ҷ.��(�Q���,���$���xbH�7�~-�aF�>W���@䚽A�V�3����?a��7(���q�%>���_]�<!U�M����A�*z�����^X̓�O��ʣ,ƦM�������ڍ3t$�����kf1�E�������Sq�I������m�IG�ɉU�=�S��u��T�H#���d![��Po������'��Tx�ŝ!UQZp�_�f9��Ǔw�T��I⟄��4�?��eű(�m�4�u��	3��V2��$�O��D��B
l�JQ��A9Y<q-k<�0�inL���LT���O��N,ce�'��[��3ٴ�?	�������X�d�<$:\���U��ti3w�C+6����O|#���O>b��g~baNV������# �yV����pl�"<���>G,�("�;|��q{�$A���v�b��)��vq�C!����D�x4r�"O� �$3��9(,�q�J
%�%�'�2"=t��?s�AXv#_t,tq�G�4@6�6�'���'��X��Y3�b�'�B��y'(� ^9$�1��*2Iz-I�$\,P�1O��P4�5�0<y��:Ak}P�ӫL�$�a��Uܓz�xѳ�$OJ����5|�1{��yb�ݘq`�O��.����)��Oz���Op����P�x�J�{e(��
���*�%4���v�
�|��lZ-~��ȹ�O'?��)�)O~�����c7@-Rtl�Dn�pr"O呀iP>Ue�%� ��G��"O�M��+��h�r��͗n�$��"O�y@���R�0!��N�d��hQ"O�� $h;������ŗ;�"OfT�rH��6�<�0�d�!��["O"�r�EM�~�*���0�Y3�"O�ȈŠW6�hm���
���r"O��(�܂<��di`�X�F�E"O�����1���ca�G��T��"OXX	�3$��R�;D1�B"O�HJ�mM�Bѣ��D�@,����"O�<J�.̥c���%��I��Ҷ"O0���)ɦXd���.�2�H��"O�T�+U��HD�D�ߚ-� �"O:y���C.A_� �p�8d��H�"O.��"<a �F�?��p"O̊'��B�(��@SP& �"O�d{ъ��#\�QB��1_�A�G"O.����O4 ��%��%P���e"O��:�l�?o^H	�DL$� p"Od�ig`��c�N�-��a"O��x�Ŵo.*HB�Ӻ
)\�W"ON%�.�@\���*�E�m
�"O����fٴ{�`���IԡK��)��"OJ¶G�+l�,��fߗ@�h�b3"O6%R��9�����dr "O� ����
�*��S�ݫ]�2�#�"Op���0b�jb��$��%�U"O��@�S�q��N��]�0"O��b�)��I�\��c ��:���"O�mQi�Һ� ��Wc��0q"O�0���j�r��F�%� \8�"Oi���M���Q%D,��r�"O�-�&�@Ht�J��Β"bH��"Oj-���՜-,i�$��,Z�ic�"Ob�˂d�{�ɀPN�>=�P�"Of� ���k��б.8+��rG"OL�aEdU#g�4`M�L���A"O�=3"�U��(x!�U! ��%{u"O�������h��T'��^��"O0�Ce��?;��J3F
@͊�SC"O�a�,o'|l��d��z�\m2�"O���aGG=�Să�,�0�P�"OX�#A��d�paC�F�'���"O�H��U-	?���'&� �R=ad"O�!0e��^!��ڮA�`�ڶ"O��b#DտY"��r�ƶ1w4�HA"O�`��B�>F�� �'�4Җ��"ONh	rE/&`dp�%���YȖ��E"Oഋ�\5�����$P�8q�%"O�<���_�q����rƄ
8�
�"O\`ɠ*�4�q��o =G���4Y��KD�C�����S�NH4d��/]�1���s�M�W�}bM�_,����(<�Z����^/��*�c�?e=!�'�D�q�̝N��9��!�|2ў��D�;UmL F����S�B��T�L --��� �Ʃ�y
� J���I�]�2�
�$5�P�b��'��u+��tDɧ��8|c�א9u,���H]���� D����,ʘl(����2�>eq��<�o��G� D��B6�q4�@�`�p��.��-1�O>�Kf-#ߘ��@O\�}\�x�&�K%__�ɑ�"%D��0���|�2x+�ɗ<;�����$ړ2����)߷���{U�U>&
d3a��.?�Ր�"O�EH ��X���c�l\$O�l��'���Ů^|�S�O����-Ǯi�v��C���a�D�r�"O��!�T'`�t���F!tJ]��\�<�U�JUla{2�E\�e@6,�4/-.)�3'����>ɳ'��v�n6�J.x��t�t �*O^�˧�G�n�!�D��N�#(�
�.E[F��i��x2�R֒�S���?��!�`�X�B�	mM����D
Iȍ���p�!�ĉ�����U9J4 �r� �!��H/��3f�P4�`:��Bu!�dA�p�Z%pR+��;]�!N$;`!��!GZ�"�
܄�āCWj[0nI!�ąt>r��@��\���(EI�<!�D�pv�槎
3��@��g��]�!��;7�TI���mҼ"d�߱1+!��S�&9���soAof���eė#!�<,���F$� .T�]A�%
�s����ē=���	�$�?f'�h�#J�.%�L��ɩq���&��JW9S�tۅ(��3zDM�7�8D�ز"k+C�����э/ḇ���ē[�^Śg�b��~R'�M�H����>cZ,� ��8�y��
���q��.ȥ77.���Z�;�����m��%�t��O�Q�W��Ȣ>�I�)E�C%lߖA�8!�f˂i����g� �M��˓��?!Q/] =��T��H�}�f1/U#Ru�ҧ�?�OV�!�L�u�x�v$�?O"0�$	�� 4e�?6��SÂ��!�J?M�&L?p� |Ib.��*W��K�8D�D�c
0~�����E�0�`�Rz��!���C�/�����O "|�D-����ռ?�k��C�8��< s�!D�,+6DƩH�F�!-Ǥ]�
�c�"�Ot��Pd�+6�m��H��-)2���[�ؘ"�"5���� ,H)
��d��=L�HC���$eIT�Q�L�`�$����E�b��e�p�K#�t��E��p?U@Q9:~�x@A�%A�x�LZ`��$;Q@C0Ŕ��嫖�g�Ym�@�I2)@�ܺ5HO'���8��$�!��4�B��Q's}l)\nfyE�(,�L���^�6)ܴg>i�q�Oʬ��/�,$p��ۖ�E��8A ��'�X�����<��Ċ+� � ��,(M�ِ����i6y�\}��Q{���s"nAy�'�$�����aܙ;p'"(�l�)�{�46ԕ�#a���sc�ЭH ���)s|��!��(aX(Նۋ0�肣,N\b ��'Y=/?Vb�)�
�)@lX{�
�l��k����4`�����G�!R!�OW!Ո���,����U�^p˅ĦO`"(��͒�M
�C��H�.�A
��-��a��6�ݕPB�H ��|�2t���b� ��FP$i��P��O�4��HDF�Ճ�5G������* @�鉃�B�bD
E5�́@l)a�0�Tƌ!g�z�SAL�-JV���
Á��p ��uD�ݠ`��?a*�����i#;��*�(E�O8�#�
(�I�T�8�!��
\f1���'R�Of�� 6+`y�1"�=H0ܳ�ꘑ>�@��'(��񆞋{��YA�NZ���*Z \�踺ろ��P�y⊜`6 q���K��y��n�0��Êe����h_�yr�[��٥�!~�s ��0��'��@s`	�K0��@t��mh�	�H��x{���*�z�(uJ��J$b���	6:$As-9����O�j�H��D(O(�S��D!���nH���%�H�	��p�a���dʶ�0�2�Oڍ������F*7M1O�����V
wͦm9��
�?���_�~�,�3��@;I��w��2^K�Ĩ�Γ>#a~�F�c�TI���$1���ʧ*3�t�9�A����L�����'�6�)��V<Q�p�;4wNT�qk�1q�,���N:E�����I�?�˓:�z���z��9��L�Ty ��="��8��[r���|~�!!ő$�� n�ŢL�H�����ć/""�R��9�a �5K�O��V��7QH(A��HVe�\�u�7�pP�VII�j�퐑�ɧ�h�s�/�e�r������mħ� �����5=�`{  ��`e�*�.I7 x�'��)7 ��afh��Ɋ��<�y�E��r�P<~R.Lx����G޴L��+��0?Y�ţqoX�h�/T�
�Đjb��E�P=s���RvB�DI������;x�.ւ%���j�I0�A���Ķ��|��B ���7&�b*s�K�bZ^��b�I=ez��T��}a�03c@�k�����?�DS�H���Ӈ� 0�Gf��a.Q��XfBR��׏� p��	CnЯ!�4���U.�� L��?��r�� &�qSQ��K@�x��b	gIaz��;�	)��\H:4�&G.�y"a{�Ґ��Y�FW�I��
B~�4MV�>���Jt�X�gƞ�}��m�����I*|-�gj"D��
,/�m���5|�VL�V�N!N*����&��io>�'DA�e�\�|��ʪiR
�݀z�
dCm�?,V40��ӧW�C�ɠ:
�� T!8�����S�2,>��K���s�g��C�c�!����a�� <#wV�z��o��(9�$�"a�0�``Фx�Q�L���ү/H�);�,�!n1�dh�<!Q�9���2�S�;:���ŬT:R�*���HX,��#��}����h9z��M@7�T
[x8;t�!	��3��$4�Nd�����WТ<9��e���A�`ݘ��l%�0��o:D����FM6i�:��B@[���X��hꑞ֝�,Rvt`Q����j�0%�ߩk�L�9�n$h�͇=?ز����	@����%ۛx�j�D�?2�9K1K(=�`m!qɚ�/������@�c�V�}C��-YL��F{�� Uc�q�X�2�$��f���'����!�" T���� !�}�L<A%C�Z�bQ��lȓh�Z5B/$�2ժ�&%hNa}����4���%a++�����Gbz	J7����F��F�@z�>!�w~�}�f��$���(��49cv!��'>:(��K��N�>8Y�#w�db૓"�hO$���ÖO��Eh���Y睇��)�U�aP�����E6�
���O%f���3P�S#rH�h��.4�T� �d����	Ҥ_�d��i���#@���)�]� 1�N>�1��y��R6"-��2�@�Z�'�	PWk	���a�dT0���9�O����;p�2� �(W)K�ry�5�L?yh��&�)@�b��t*�uX���0c�
�|b�$N�o��A'O
L��\��h����"cA9d��=�
}�U�7`��Ro 9���0K�Ό8�:$�0�`����%a��"#R\����M��Fyb��\m�e�
�b�R]���r�ճҠz�NQg��O��X�,<�O�p5�H�>�u���ES<�"J
�\pQ��&WV?�b�H6�`���Kv9����߂i��D!W�I8�ԕ'���g����\Y�32ɐ��d��@���H֦��-��	�$��1E�r4���p�H�g�	8R��j���!>`LCH�6|���c� �2���B�j�h��H�c	�F���%�r�PL��E��:� ��/cSZ�B� :�8D�L:?�#0�&@�t�ϠH�n��G�����Ae�L�,���15^	�I�
2F	���N�gF�<W�0 D�`�`�����	e�$�PEn�A���K�Ę��y�L�Y�>t��ڔ.e*	�f"���0?q��X/'��ɀ1�N&#>=���).
��Ϝa?Yq�H�	XP�Ԩ��<f�b/��Q���P��O�JX��O�x6��Y�����Ըq1�|r%�'}y���E%ƌ���An=�H#p���y�n�=��X"���)*)�5 �E�gh&���
�'BJ���8�A9ܵ���ͱb���S��
��ɤO�X��*�E���5 ��v�v�;R�������X�\�N�(]e��"?Z���D>z��	����'U^a�		mT� �o%ƈ�J��ʻ8`��J<��nM�w񱟛�g?�@�ó(����&��L�TS�{�<AwC�FL���
B�pC���<It�ǉ���� �p˓H�V�<9�CPj�*l��bʵ3~4�LQ�<!e�͵^3PUXe,̲6a0��䡋N�<�g���� ��U2��8P�ft�<�����=ݎ�K��ݲ#�ÁKNs�<�/zW��a���&�!���@G�<qC��1r���"��x�<;$ IA�<�҇.g�x<� e7�%Y���s�<�ƨ-AWf��ȳAdP(2r�v�<)��]d���b�.z�}P� D{�<q���Y����	��:�������w�<9r�	����&M�(j�E�2"Fq�<)q��d����O�
z�� �j�<P+I�;p��2a�5��m{s!�c�<Aca(h��@�3���#u(�;R��\�<��b\�	8D��V/}�� ��X�<���<xF�x�#,eb����Pl�<� L��b�O#qG �q�$qɄ\S�"O^Iz2]\x�˕NJ��|"O��+U"]1^�j��p��,Q���1"O��(W(��
�s�熾p"O��4I��F�0l�VFĳ8x�-ۇ"O,�[q���(��h¿1mi�G"OЈ{����p�ㆤS�0��x�"O�eY�i��/���dd��q;�"O���@8���雄;��3�"O�D ���kې)b���Ua�"O�=拕9��(�d��3�1�U"O�D����"?� 42�囹>P�ԋ�"O���g��H��/'BDxq"Oh<�1�E�7aD�Kb��5Z��"O�H�d�6"m�9�󨏾'��7"O���D9[9�$�!��g��Y�"O�H��*��A6$����
1���C"O&�`M�>s~T�3
��Ԙ�a"O��3"�**S�a�S=y�i�"O��2��D����Y�hЗ"O��� o�;�,Hr$�ӷp��Y�"O�}dG�|{�qC�%�
E��ĩ"O�p�-�'&����G`�L��"OF�K���4��1�5�N�i��W"O��DEdTܰ�!�	p�,X�"O"52ͲZ:!!Qc\&�lP��"Ov��Bܮ7�|������&E�e"Oj��D#����8��L�`�ָS""Ol�8 	�7�a`Lܾ
��Q�"O~�!�W.�5��L�}l�}r"Oڽjk�V����OJ�=O�mSG"O���d<^���N��D9��j�"O]���}�N���,�34$�ʢ"O����$gn�1`1-|!pDk�"OH�DL�2��":&�Mc"O �K1��^{4�qP"�9M|-p�"OT�����)_n�8C!g�H!�"O�ԉD��(f@�m"Do��&D@hF"O��rj;-�P�8r��P�*�"Oj���dQ��`���cR6��"OFd	�3�� �H0.�$"O9A̑/
���s�]9�<���"O6pc��	A@�Gc�6�0@�w"O���.�	����\�o��Y{�"O��1��C;y��AAT�41ԤH1"O�����p,DhP*�Hh"O��bbo&д�ط�T�R���"O�ģ����Z�k �lM��[#"Oܘ`�@4]�Hѷ�H/��a"O�{�뉷s8�@G<58ʭ)�"O��s&�N��%�Z�Uh��2"Oֵ�7�T�-b�ѰG(O�4�"Ot=�#�
*����2�pd;�"OB*�* G�y��E�+�Ḅ$"O���p��$oȈ,�퀲=��Ѱ"O%���\�u��-��r���"O�qٷ���d�ݑ���%+=�"O&��MF�J��4��d$*ؼ9w"On|Y2M�12iX���	_8��"O�]a��I�D�(�ڕ`�O C�"O)����7s��Y���'Sf\�Y "O��"��بk����.�1d*�RE"O���CK�%@B���%��<nH�*"O*�c��� I��ڹrT�4P�"O� ���`��k3�e�a˅6I�=Rv"O�d;c�\�v�ɸ�*LN@R���"O
�A�
�4�:�ӲG�h�~A�"O ��- ��]�'��٢`"O
�B����ʈ3Fk�29��"O�M�a[w��R7'Ĺb[�%�g"O�"���+�~	��k˄ 鎵k"OX`� �2kF,a��Y�7��4K�"O�8�$��a�����)�*}bf"OLc$�V+�|��i�Ns�""O�D9 H�=�*�!�gS�Po�X��"O�a���\�K�lI2a�ɨS`�K""O� 0!��MGܴ*�#Ȫ:Ѯy  "O�`Q�ߔq�j��D�j�la��"O�=���`��%Y��T0�>�#C"O��/��7^L���Č^Քs�"O�<���I�9C�d[�V=�a�4|O��a�'N�a��$B�Ã�JČT1"O��	�-�.������_���i$"O�Pkb��p�r�������!�e"OZ4��M^�z���ܤnV��'��U�ÐS�Z0��
F$x��' ���4(�=_'�]�6��Wպ�'�����h�5o���f�;q���'�� RU�	b� 5�%6U��
�'���C��/7�H0$탻-\��O��=E�t0Ra�㊝B�E�fM���yŋ-ʢ�����>q��M%�yb�� ���p J�b����BЮ�y�E	�do4�{B��<S�8�Q� )�y����5ȘD;�%X�Gc0y揙��y(D?s�����O�"?^��ȴ��y�呁'f�0-�"Y(Y�-X��y�_.ƹ�䢇%hB~�ce�Ʌ�y2��g�(�QȒ�Y��]�4L�yR�8t�
܈unYn�|��X��yҭ�+�����,P#�`����C�y���01|�	��X
���4���y�BZ�_Z��x�.T���S���Z��C�ɞ
9�G`���)b`�4k�C�9#R8ꂭ�[v��描�F�C�ɪ/N��@�5ej�IV�Lc-�C�ɀe���D�/+:���CM.ͮC䉏
�h �Bٕ%�x��+?�C�(PB���ҾH�f�Z�N�"YnC�?7{�u�ω08�zQ-�3>�TC�I4?��0qdE2SSL�Q&0%X�C�Ɇj�l� ��~�:�ѯ'��B�	�fNL�"�'#pH�R�,S�bB��P��#�$R'}�"4�&gZ?((8��$���&�@����(5ih�0�G�3���{3�>D�@9�C��3ƥ�v��R��X0D�Hb�`M�op���L� fId`��	"D���N�1eZ`w��9!�: ���!D�00�V7(p�4=�8d���$D�HP$MK%_h!8��C9%� �c�'D���_9�T�1MC�WWֽ��%D����%^<N�6�T�@!o|��)�d$D�b���5@9I���@S�(u�#D��s�J�	$� �h�5�>EH�b D� �u�Z'N�p���8Kuv-CA�>D���4#M�G(ꤹ3�?6�B�(�:D����F��2q��` �ˆ*2)*�n+D�h�d�@��@�05�N�mG-����O��=9��� � vX�0��}Y�hY�e��$i��z�"Ol�j��(M�&�
�eZ���FQ��o�w�'�Q�D�1�U���q�N����� D�T���N�D{B����#sTtl0fK;D�(SCH��!ɮ�9��^?��x�C<D�����R49��0c���)'�'D�@;3��?���{P��� ��1'D��DN�"��{e�֢p�P �:D��� ��*���ؠ�< ��`@3�y�x�=E�ܴ'r�9�taǈGg T�� ��E/��ȓk���$���@G*�<)����q=�������>O�08գ��Md���ȓ_�1�0$r�[��ߕ-آ���X�R�
�CE3z���S��YADY��9�䐣���)�2as��	^����ȓxJ��j��T+kXB�h�f�3pXa�ȓ$��2�H$ 0T��2���ȓzLi×F�x~bt`��^G����ȓY� 1i�&F��eL����=��2��H��Vd�0�@Q�D�d̐U!�^k�.�����-�n��a3J!���X&��V�I z��p��ՕI3!�(uՖ Y��V�;������!���''.��IU�� ���4v!�D ?_*�qV'�9����P LJ��=��w�J�K�oYJ5���پ0D�=��iyb��D��B�]̸`g��\�(��3D�l	r/�/n��ivㆪbn��'1�IC��	'�R��r�
w�Ɯ/ʶ`&9D��D��U$���Śl�����y���%kbAʩO�gܓ�ļs�;4 T�M|^~M�ȓw,�B�杋?�j䱔�т%,R(1�'\�	)7ꕫ}4 ��!Z	*��C�O>�=E���	j�$T[1,G=[�v@�2�B��y���|qŭ��O�P�WJ"�y���:�d�@Ԍv����lN��0?�-O�`���@�w��cD�u�,�k"O0 �NB9/`UʐK�M�$es&"O�1XT�
1��,z��� "O�l��L	���=Bg(� q�:)жW��E{����8G��!�7�G�?x��a�J\b!�d�
��7 �+Np�
��ۅsa!�DH4l��4��+B�B�%ڋZ�!��ּ��]�P�V+{�ӳ�R6@��O�=%>%a"$"-^�!���X���0�8D����e����E:�'� CW��r6�6D���u%�al���ű-�Hq���.D�X�`I�Kt��℁7{iv�ڧ..D�qF�ǳR�reSM��!�hz�)8D�����/~�4qa�30iB��!D���a�pr����ݧf�0��e D��1G�`P��j�$u��k��=D��q���~E�[��U�"p^p#)6D�pr6�����P�@ �ɖO/D��	��AL�}�+�5"���+-D�j�I�'�\p:�`C�:���1�.D�8�Iʨz]�L:`c�
z��C9D��3P��8���"�Ȝ�ݢ��8D����0A��`��#޶%x��#D����HԜs^p��F/؟��H�c�4D�p�r�/�	C�%W/�a�%D���`��>|-��#�lOZ��-0�0D��(D�^�[^����5>��̢�� D����z�H�	L�R�Tt�SJ+D�� j�qᏒ�D|hAǦ��K�� �"O
d0Ae�-`L�	$�V� ��P�"O��v��5d�*���ʉ3N�L]��"ON�Q�̵n���*	Wv�V�B�"O�\k�Ɠ0���r����4"O��&%+J��]X F��lU�E"O��ᦋM�Ѷ��D�L��"O04�d�׬Y�v�x��֦`�TK�"O8h�g�60��:�	�dd���S"Ozaq�.M�N��8��i_�&� cb"O�л�<]�A�pI��a�t"OƱ+Q�T+7�I��N��0� E��"O����V�{@q9 �Y�a�����"O�Q� ��A6*�������W"O�4C�G�5S�jB���M���"O"L�j[�G��gL�5�E�B"O��Uh�O` ��J�E"O�QQϒpP�����O�z�""O*l�7#��@5�b�cƂ��E"O�����	f
4$CeȸuT��u"O��a��-b��� �E�-A��(�"O41��'�5~��0���iQP�jf"O�yxV�P t�С��jnpT!"Onl�p���&�dh�2DH�wT9��"O�P��@ج�+"���B� ��"O�y��B��2�� �;f�Pa��"O���c��t��ӆ�WnĠ��6"Ot�b.v�i: �����"O�h� ���;b �r�]#�y��ɥZ4tubd��t�C
�yR	�8�z���3QUB9�i�yB�C�^6�[ĭ��쬱���y2Q� �X��	�KR�Rr���yb@�#:�A��xt\]�@�\�y"�
�xU�M�b���%$x�1�dP�y����V<�|R0L��uc�Kי�yb��iLl:%��,] ������y�ʔ����J�g<,!E�y��PtW��b�șf���p��#�y�靗gi �ԃ�,`%�AYY�C�I_���c�F�;�J��-�,/*�C��&`Ϧ�{��Za*&�*DC�	6@�T��� 'KV��hP�.
�B��--����2z�JYB(N�\tC䉲瀑��'ّu�d8�k�*(:^C�	i��aG�Q�w�P�!��ʩt��C��~��4�!�����+�ᓴ!u�C�	?{��mZ'�1VIJ4`c-�?J$B䉇*yz����3�:�ːa̗:&�C�s̴X�э E2T!�T�c�C�	�[��#ԀX��l�#"�R�4��C�'+C�X�w��~�`�i^=�xC�	(
� R�ݫCoj*5��A~B��!%k8m��'�.t@X�b�!3jB�ɻLZ��/�c$+��i+&q	�'͋�B�-�-��FN�aF����'�b�e"��t����ce��	�' ,!!�*�
���rJ�`��ԡ
�'9�<H�Ǖ4FN��M�opH�	�'����6���*��F	��`%N)j�'�&�B�"]oe*�S6'ӆ,]���
�'\��VgS�#�Hd�Ɔ�Y� 	�'���SH�V�����G��պ	�'�H���g@4Cx����=B����� &� A�={��`��F�F� a�"O����P5,��A4ˉ�A8�Z�"Od)V��(Ip�'*���-*�"O��2��"RI�Ai�(�$�A"O�d�B,�& ��ST'�?(k�H@�"O�$�6�W�7�}ѥ�b܄�"O�铰G	�[0U�&
�yܡ#"O`<�&�_�O E9��M�x����"O���!K@@ i���Ih�x��"O�5l^�+rHܳ���S&9i"On��V慜Z���D>-k2ѢT"O"Ɂ��}q�T��0=��@G"O`p�#gA�$U!�Rm�91�NUz�"Or�	V�K=@��� ��	Z���p!"Ox)z2I�b�`8��lK�bPh �"O���"���42W�ܺ2��x�Q"O�(S��Pw��JًI�(��"O:\�gĉ'(�@���ɕ�< "O��Em؄(R�b���)D�����"O
uB$D�B�J÷oѤND�s�"Ob@�F��&v����-M�X��	)�"O0�K�I�t� �a2J 9�H��"O�$�%�ͩF��x�L����0�"O3��X�
ٮ�z����,�AS"OBT"b�`�A��� �,}��"O�˂�ߖ�PԻ�86�I��"O<D�1��Z��5�\b���un�+�y��հ�h6���������y2��*G��A��a�)�B���Þ�ybn֛*��RǞ��M�e�	��yB�ȕx�$�t�� 6�,�S��;�y*�%�hŘ��ȋD2^����y�['�8#Q�"D���3���)�yb�('F�9Z�H6MSZ90Ũ��y�LL&�t��F�9���
5"�	�y�(PT,�A�q�AGK0�g���yoL�Bb�	�1�V�P
@�fF��yB%]�Y8� �-�5�h��L��y£�\+���"�!V��[�KC:�y�,E�U��`�Q�T!b�+��/>�ȓP�Eڗ���v���R'*�	m91�ȓW�)�@��A�Ѩv�C\f�ȓn3ޜ8�CSU��)���sD$�ȓ��PZŇSoD��w��=^:�H��+��{C��咀��-F�~�;� !D���۴w�\)B��� �I��;D��Ag�Ն7��� BC=}�fm��,D�S5˔E�@����!�*ݫE�%D����W"H�� 
 �K5*�B"D� b�A�y��"�Ɋ^�ae�>D��{A�K�F��u!c�H-L�Td�">D�T��ð@2h���BJxQ��?D�<���Ib�m%2�	D�;D��rnE�wM�h�R�1WkN���C8D���$R"~���B�=��rE�5D�ܠ�* Z��� �;�!C�
4D�0���1B�>�9��'.���DG%D�(bCbV _H ���N����g,>D��!���
������X#R�����8D����mD��)r��1"�qؑ!6D�4s�FY�2޾�פW�����1D�����h������%@�<B�	�}��0W���.����A��DB��}�J)ygc� &����i���B�)� ����F�t_8�hn���X x!"O�1�3M�x}h�nQ�lӲp1`"OPI��KS̉�ă�t�>-��"OT����5	��<�ǩ��(� ��w"O8�z�ԏo�����&��.+h!z�"O
�f� H�sG�	�+��h�"OXq���ʌT%^LpԇH ڊUR�"O�HQULŏb�>qq�J�M�``�"OacS�նi��ъ��ԕ'��S"OH}�GQ2�`�z�ؠ8
�15"O�a!k�|�0�E��x+^��"O��Z ���*�P5�<%�Hk�"Oz�� �S���b���;�|[�"Oz�!� H�����ꁀ.F�{�"O�e��j0��A-tX���"Op�*Q'"Ј�Ӓh�gf�Y�"O lR$f�Lw��kr��9Lg���"O-�ũ�1Ft1���H%W/�i{�"Oj����'�R����Wr��u"O�������R�qt�Ŏ'T"P�"O��,�'��d��nɟb���C"O�%��oą����@ �U"<J2"O��B�lb�LM����B �I�"O8��$`���9�M�
y��1�a"OR�A�*5���e#Y4K�>%�"O�f�� a�u�G$^v��@�"O&���GF!���ȰbܿVEf�2"O�٢�(�7@�d
�+F�1�= �"Ov�Qb�K�B�AՓh�
"OЀ�тK���1"�%\ �!yc"O|$�W������G��~�v9�'����SX�a����3Kzv	s�'
�e`C�ɽRV�������p��V�Z�VC�	��d��դA1B�ʥƙ7@lpB�I�{��A�+Wv����V��pB��"[	tB�n7F,i�-�8�8B�Ƀ/�0y2'�!X��T��k�B�	�x����g�3U�QX���#��C䉽`��Y�7#ܣ ���3b
�PzB�(�L�A�^�/�~<�w�,qp�B䉘<T8؈w#.lC���H�~��B�I� �\���@ ��)c��5�B�	���S2	��]��#1��z<C�ɼxH3��@/x:��3�R��C��\ �Ѧ"�"�8���:l��d"�� ���+ՠ��M��q��e�6�5D����B�l��1k@�K$R>� 5D�P9/M)5+�DPN�$p��5�o3D���ξ`�b����1'���۵N2D�й� �%��i�p`��UL�Y�/D��j��΀P*d�R���86"�-/�Or�4%cTp��g^�s!r��ƍ!���<�	��0�� = �c��OB�B�	�4TZD��c�'d�^8�C-S�7�B�"lf,��i»J�4��3�� `SlB�	9"9�X0�\�v[\�@��Q�K�8B�I6 [� @`l��/�L1@Wڙ_�C�ɔ<nt�Jw�ש[�.i o�6;�B�I7K����5c֠n?�K��(lC�ILD���b,#sP0���Ş6e#`C�Ia���Cp�L# <%���ڛ]�P��0?QҢ�:]*t���q��a"X`�<!��Ċm`2*"č5}�ZU[4�_�<�CD(��Vfۊ%� ���Wa�<� �e����N�ذ9� q�`�H�O�tp�oܚx,#��ׂ$DqQ�>���D"�&=�x���[��̢䏛H?> ��
�H�ju��-0N 횁K��E~lY�'�0 ��N��Dr�k	�Bz�%��'���A���+:�ph��,zV���'�e� ��7	�S�k0IV4x�'����ͩh��l��E��~cj4��'
����A#m @(�%ݏp����'ΌyH�J�������eV@Y�'���B O�z6�є�V�Z��Y��'E���QȎ�R/9i�FM�Q�x�	�'NV�gG����v	>�6ى�'��L*��+rBY)q'P3$�HA��'Ah��KB�I7x���\"
�ɘ�'bz��6�*j����q�.	Ȃ�����$.��S�qeja1�Ă�7� Pb�F+6��pغ#ev\рA�!V�Z|�ȓ  ���P���)1XL��K�cW��ȓIS�ʷ�	�n��0ᇆ�hv�ȓ<��0S��u�F�R��r�L��ȓe������:���T��7�����X�P|j�Q�~��l��ދ'`¹�� ��;F��N�8�fJ@�Z��m��L`�I�����]#��.Z� ��ȓ�亡l	'���
T,�-��l��^綬r���9��u�Gm
-G&�ȓ7�!�\�߀嚔ϑ)f��	�ȓD4\�u�ڜ:�.! &O���6Ʌ�Ns�r����g]�I��g�h���2�4A���̝*T�=I!�K+m9����/9D�+B�J�$�^9QUo@�e��]�'Ha~"kM1�x�6��k���T!L��y��Aʼ�� �65Z��t*���yb�*"-�]��O�~�0��=�yr�B�K��L�'�G�{x�I1V�ǘ�yr�W�b�RnY&82)B�&�8�yb��C
���OK�;����W �yB�ƛ_�8��'�H5mE����$��'k��OM�<Z箞�q�蓀 �<*��
�'��y�p!A�=�,0Ю�?)�
�'�"2VC�$�(���7���'�8��a�6���A���q�.���':�H��(LN�l��D�f'���'���"j�N9n�8�d:Y����'Vj�s$�^c����h��S��u��b\�XD�d��61��a�h�;sVJ�S!A�y(���Xd)��5���`����y��2D�J��:d�Hy7���y�,Vtĥ�3DX�Q5�&
�$��x�J�&dҭs�f�g�D�vkB�!���;V��(v�Y�	6M��ʱZ�!�\	<��$n�c���#`	4��O����O�"~B���j B�Ȟ�
Jx��n�a�<!��uZR}cc��#TD1�kZR�<��
�N�j�T-_�x�eeC�<��-�.EB:�hq�
��� �Q�\~�<A዇,�V���'����
z�<�T�	�\Q�E���D� �c *Ry��'�A�%Q�V�=s��1s��X��'|l;��O6�dcm]�A!�0��'MBQz�\�C�F�)a!�2K>X���')�P!���W���0�ШQ&G��ybc3m�`i"��V�|��(ѫ�y
� �d9%�^�8�f�!ү�~x�5a�'�!�DՇ6Tl �IF*�n(4%�F4�yb�	�I���1�;+,�PKǊ;oX�=���}��( �a������.��q�ȓ.	H9P �U�3,z�s�k[([���ȓ�	�Ѻ�>��#�Ɋ�e�ȓ�9]%�N�����Bj찄ȓa ]ء���o����H��2q~�'�G{"�C�t-T2gܤڸt(��M��!��A�}�����+a�d6�^x�!�D���ɐȅ� MH�e�W�!��UtHb���ϫ6�V��$@�Z�!�d�㆙8ӊҶM��|
d�ͥ8�!����Hr�(�&d�\��+ 7�!��F?x$�Sf�ϸL��R�'�n�!��k�� L�9��2G���!��ؤ=�)��MR#L'��{-�!X��Ol�=���%��ܦB`~qxU(E,H%2M)#"O:�`�ٻ>w�p�& ��"`Q"O�)��7C����6>��p�"O������BV���#�4Q���E"O�c���8zfҴ�$~�2"Oѹ4��pA�г��?Ws��	r"O��q�/Zy�x��-�=De��|��)��;|c��3���2+:�@���^#(C�I�xU,d��GͺM�`���ϣ"0C�ɕP�����LD����3B�:c"B�Ʌ#*�Sہ`iVAP�K3u�C��a�Ǣ<fā@o	<�C�ɪnd�Ak�R��	�d�>+�NC�	
ڸ<k�e/e��TH�C�I�Q?����ԡ� �T%�h�xC�	���h�@��
[G|��g��<�dC䉺=�h��Q���
xħӖx�.C�ɞ7���գ]���	��b�LC䉾(KV,���wf�e;t�C�I1 G\,Jg �u�X�A�� �B�ɿe�tyE+K%i₀���,7�x�H��ɵ�lE��/�9q$D�d�,?�B�	]��Ǝ���r9�1,ۦ��C�.kTڢC�L�(�I��z�C�	>oJެi1���V$Fu����8�'��qɁ-R 9;�o ���-O"�=Q����?Q/��ԆAl�ʍ�s)
�!�ń]�B	c�Cݐ	�jT���:J�!�Dжִ��$J|s���Vd���!�D�:^զC�Ȃ�v��\2���Aq!�đ�$L�G��'���q���l!�$F("yA��F���&��T!�%3:|��p
�sܮ�S�/'I�}"����J�Q"�8�Q��:i�H�q2D��3fư1��������p�=D�+�JC+ ~��) ?~�IB��;D���s�ΓZ>����r�M��8D����	X�`q6��<5x���9D��C���{�q�%FD�n"nIz��"D��@�H�)vZa�a'I6����?D�0��tTz3nC�9d�<D�4��9�¹��
�r~`���i-D�0J�·>.f0�!�`� � H��?D��+��V��4���Ηs��a�u�<D���#:iC
0��(
)��5�o:D��*"�A<o����`��;ޠ��Ս%D��A��E�GH2IBG�P�=w��:�%�O��S�? �X:�X�#�:�ۄ���E��L��"O��2�G�x�^P���+A�̱H��	}�O���;W��T�.4ಆ�)�<���'�
9��� h�6���NÕS��i�'�A8��	��T!�(PCR��'ߒX����$PF4���B���'>V����;�L�(���(.�(��'�P(;@�#����£"�VU��'���0nX�B��гB�R��I�'bzm�B [��(G+�.9��E�����$!HJ��D�ۖ5�Bq��ӈ��a�Խ;�L����7K����ȓ~�x�g�u�T��rN[�x цȓ|�f�ÖE!d�I�Ǣ �?��U��b���� ��%�R�����:읅ȓfD����˽3c �f=2�<���G���h���ܑ��mK��R�cgm_C!�D� V�j8���Ȕ%Y����4!���gT�A��N���Qfe�w!���"���9׀� ���W��a�!��}p��sO^-88"�K�)Q��l��8���>J	�Swn�4
y"2N3D��k� �l �#Ȅ6��`�-D���R��9&���:t��X�i�!�*D�dp�H���}RF+��\|�z�g'D���	�!G'd�H�-�v<P��D D���eL%]�v}�$G�e<q��E9D��c�GB
[
��seĂ�ntv�9c��O��=E�$!_O�������L���3�M�&(!��9�pr�/R���{�!�y�ɨu{@`���ۅZ&6�Ҡ���B�I�0�0��rŜrzTe�`}bC�I�>t��笏�L6"�w'��}�DC�Ɏa�H�:$��n+��3���+��B�=9;
=�w,	�3Lx8���_����0?�4.��<>vec��(a��Eڤ`KX�<��H�>�*��È�29n`2+�M�<1�bA� ������&v��$�օCK�<ࢂ,-i}H�e���L4�'%o�<����~o��y��Kf�����l�<AF�G�.`v��c�z���B}�<1��&H/��CK	mWh�a��y�<q��V;j��̹���:��q���r�<iD# �.!F��1)ٚqb,l���y�<��(����i@�5�$A�p�t�<����J�,"���e�h���&�m�<�P�Ȥ"UV��d"�KZ2���iM^�<���ӑk����O�`T$ �͐r�<	���9~�y k��/H���Q��o�<���C�'w�Y�ٔOuu�NC�<1��߽
�K��C�[��:�A�IE���O�	�C
ϔ[xZ"��';W@�b
�'l���Xh�f�r�8m���
�'8���jX�En�x(�D&|��2
�'ʀ�(��$#�d�3Č~E
�'[�$R�m@�mn�$�R&N/G��\"��hO?)f�܈0l�T�Ff��\���NA�<�@�R
�(u 2KʁP8����}�<ɦÐ%!P�q"e:*���c�Q�<��CĔ�0�Y4Ռ DMZV�<�P�D�t{�<��Z) U0�a�O�<�SKͷ@��`��\'rv�j�*�N�<��NBE3B�1�	I!h@,P�i�G�<��G�m�V�ٟqw �۴f\E�<� ^t)2�ӐO�M ��Ĵٖ�	"O�$���#/Fr�0 �E`�L��"O^L@TDW�N����1KJi���IG"O�a��.Uc @p�c̡:�š�"O�DK�N��>��YF��F��P�"O\�jG&Q�,c���$���jS�'Dў"~"�h�ڲa��ϫg��0��옗�y�*Z�H��镸\�������y�n�%Î� 4�+b�q	�yrG�E������( 0���+��y�E�>Pxrr�D$�)*֩��yrn݋�9���q�b咄n��yRȗ�
JU0%^-h�>�)�O��?	���S�L76(�¡FƵ�6�
�)���ȓ)I���7#�A?���"��~(���ȓs�ֹ����U*ݺV
�I|e�ȓc� ,��+!�T#�G�[J�5�ȓi�x͔�`�Ā�'�M!RM\h�ȓC5�R�KXi:�IC � }UF���(�PL�9 Ƚba��J�ܐ��k��J��ډ=��lZ��4p���!�20pv�Á60���Gl�L(D�ȓRT���,�*Ֆ�b���	Wh��c�m�1�׳T�A���݅%#8Ѕ�c^
=(��n�Q�EC�!�����J��`;��tŞ9�m� Mڞ}�ȓQ��l�fԈ^d\2� ��}�ą�q�H91ЪU1W��X��E��l���B��EJV#Yp�͚`EǽN��i�ȓqg,x��\z���QAnǓt�l��\���KV��)-�����69�$��ȓ�2O�/��qs�10�0���_҂�86eL�>�:�J�hV	.`��*PHx�F#-#�C��#��p�ȓ8h��xɤm��̻´8��IvZ����<4�����ʅ�Y��1��:����>}d�����G�T��tq���
�0������=b�9��#;�찶��+38j��&�2Al�5��2�<���c�)xI���\(���i�N�<���0$D.z6G��r���M�<���y�Y�3 ˫a^VIbs	VO�<)6�R�@��B�d�[Ol� �I�<�!N�L�
4��(�J=U6�E\�<��b�'�.�!�*]��x r@�<��Ǎ oi���R�"���BTJ�`�<	��ްش�����t8&�`F�Z�<i���'d���&��pw�) w�W}�<�Ȇ ߔ���t;�D0%�LC�<qTK�\ۮ`*j\P�E�� �~�<�6DŘt�a���X�سQ��Q�<)Ұw�J��ĈqXL����s�<��5 ֈ(��,�03h��m�k�<I!B݉u��C!̀5ݎC�H�d�<!v��13�yA�D�x�p���Rc�<�a&��,�x�Kd�ܷ�� ����_�<�u 	�	�1C`1mN���@\B�<�'�_�h�2���A,uR���I�{�<IW,өT��$�b/��=����R�<�q
Kn,,�Xc��7r]��O�R�<��Gûj5�����?����S��K�<yU+'l�IbU@ՠ'o�U���BG�<�7��N��0�0n��d��B`��E�<)${;�X�S���7��9) ��f�<� �L���_�����kVLi�  "O�1��ȕy�j�2�_mPr�Ҁ"O.���.�T��}�UF�=zJ ��"O�Q�͐�f�2��N�O8d�ڶ"OT��m�T}���%5w�>�"�"O&i���<E:8��,R�<UdA�"O�iB�kL���!�t��5� ]�E�|��'�azRkÑt���0+�.�M��-V�|�!�䃩����W��'t��q�֕Y�!򤍰�|z�ݍm����G�=i`!�$P�*���*[4@��#�K!D!��9z���ڣFV|����$)!�Ā>R��0�!$ Ѱ�����/g!�A]�L���%ׁD����o���'��	k���s��D����P2XD�)`B3D���C��6n@ޑb��[�a&�e�Tl=D��Qu�P!?��q )�(�Z�(�(;D��AR���^�F$�R�X=�:��	=D��y�IEz�����2C����=D�$�'L34plI9�Z�d8�p �6D�IqN�,#�0�f�XEd@)�5�	s������S�N�5�Fev~j���@ D��bM�}�89 �ʇpdj�QE<D��0�� CP��C�y����(&D�	��F�&5"�{��܇	��+!D�p[u��01V"`1�F&t]� �g)!D�(��n��'����.��^�T�:�=D����)�6�X��Q)�/D��ڦ9HUs"�r��9���.D��Z���ҋE�x-���I*��B�I�,@�0DNɻa,Y*%#	�w�~C�ɕt� �2��u�U�Cn�!�jC䉪Z���㤇��W����#��B�>C����X���K� q&�N�RC�	\�!����i�j(c�H�z_BC䉡���ʷ⒫z{F�a&P��C�#u��E��Ğ�V;� z���	
p>B�Iu���;d
��V�4��`^�0R"��D4?q5ʇ_�8��m��'��������E{��郉
�|}�3��s������ ?ӲC�	��`�EWE+�ȱ��VפC�	4Y!ވB�ܱ��<0�É��LB�%a
$qaEA�QЪӢ��I$B�	�l�C&*�L*� �C�Yo�C��-X��a����q���*��Ƅ3�����%?aV㐡W��jF%H=�`<�a��\�<Ѳˎ�4������js* �wMs�<��,o� ���]�|5��Zd�<��'I�X:�aGN֖l��2FM
U�<!�c�,O�hbs�-+��q�a&�j�<���ч!��,�Ӄ�*X��`Zj��<1��\�4��@���"��]��f�<��L���ҥ�A�(�D�Q�KΟG{��I�;?�1
�I�av�	��I8�@B�	7c,��r�������'	�yB�
~����iZ�w	�l� c$<C�v��!�S�W�.QΙ���FF^C�	IB5�Ŷ
�%a�iES�C�6 j�)!'{��I t�^�lt�C�Ɂ9���P�	)l|I����:ܜC�ɗu��!$䂣vmr�)5�N\3�B��$X�8�ID�"A ����L!?��B�	�QY4�hr#��T�%��.��#urB�ɉn�,q�s��\�*�!����B�)� R!���w_^�! ��kad��"O�I곫@�[+��N޶?�)�"O�e �H���+g��Ec���Q��F{��Iʫgi���L
����^�K!��	'���b�y�.��b �S�!�Ėr	H���I�`�V�  "C�!��Z?�`iP���1�p������`!��3\��Q*'��3�� An�QG!�DI3;_z��`m�X� `mZ�.!�$ϗ%��]�Fa�^yT(Z�ʈ<*!���6�U�$������+Y�3�!�$ǣn�$�2�IG�X���T�@�!�d/o�&H����v֪�"��U,i�!��.���B�ٳHq mj � <8�!�Ă�+�z]�� cK0���&{�!�d@�NPqt�N�]B��
�!���=�\�!U�$0�,�Q?*8!�����P���'��#��VFG!�DF6p���G�ֶe�3�ë/!�d� �Nq1#&�e�.d+aj��M)!�D r�������}��� ��غ !�dM�&?��c����S�?�!��^N ���Erk�؛��|qџ�E�T�Or �[1���>�6���,į�y���>��(�\�7.6P����y�h4)�TXVW�x�Mp��Y'�y��y�b��o;�h)�
��yD\ P��R��1k��2���y���n�����m$�)��L��'ad|�эT0o� �ІB8_`E�	�'Dfeeð#���v���ұ���hO?���d�7#�p�r���c��V�
K!򤝐ndJx���Q�M���Y���y��	�<�i�Ňp�0A�'*D�t�VC��e�����=�Luß,�.C�I�1Z �����J�U�� ~l�Y�'��d��B=b�T��Qȅ�e�b}�	�'�&� ��K42�xѷG�=S"��0�'�!���;o�pq �70�V����L6!�$�8�a��
AU���/�?%�!��xI^�cB��,}L����K�!�$��!�!��%I���AĀ.G�!���"L<lY�2.�Z���lA�
c!�ĉ�Y������o�� �Ub��=Q!�$�x>l��r$�y��Sg �1HG!��Z�]���Sr�رlZ���`ɓ19!�:�u@��J$ƽ)�.�u�!�dG�Za�	�W�`1�V�s!!�D}���r�#��q*V&S!�D����-Y�r!���YB�ѱq"O.T�@�і0p����<dF(�w"O�U�"לD����?)�ӄ"O8L#�l٢#��t��_qG&��"O:)�&�?.aA�*-޼4�$"O�D��,$lz!� Σ-!��J�"O�q�M�7����B`L�b��1"OR��
&H��d2�-�9\�
ݱ�"O@�I#E������U�HV����"O~5��[�S`.�"/��S#"OT�`���O��Hh��3>��x�"O.���y&�h4�O�S��{�"O��(�#%6@��A�V�U@8�"O�xb� {���K�&�BEX�"O䠚���,����*@��"O� �h�R�"8f%x1 3@r��`O��s6,����	A�#}�b�/D� ��N� K�$��Ŝ�Pb����@,D��C
�@�H��h��yꪤ�c$7D���2�f�Xz���,8���sP�4D�`�#gɼ�r$���ю,��bl1D����&΂~��ȘV�̧<���b�.D����2Z��S㋆&v���֩2D��x�E_��5��n�L3X!@aF>D�H����<�i���N�ء��&D��	v-�$W^����i�)�
��$/D��P�nԵn�"�)�B�hJ�c*D�Dd"�o���@��?���=D���#�m��M���O�b��ڷ�(D�T@ �$)� �!/?$���J"""D���'��n�nPꇢ�X�@ђM2D�A0m�H�XP�3U8���$=dC䉗���y���x�T�ر�N�	
C�<6X����5`rM	��B��B��+O�}k����R�,�sW�uxvB�	-RbD��i��K��1�tl��F@�C��Gf4�X�nQT��bg�Ǒ!��C�(?ψT B`Q��NHE�BB�ɖX�l�v&�^�И�òi��B�I�v�J0r!�Ӆw�n�{7���gy�B�I#����B���z���Bü0j�B�	�|�⁁�a�(��J��AX
�C�I�M8��i�. bH��2��`R�C��=i��"ň�3$H#��6��C� C`)[��G�k�8"㡟:F��C䉘E�L]Y�f�5M�F����\�\%4B�ɊH�`(a��D��,))E��c�����O���q��IQ$�.*�Ѱ2*[�����#>D�4��(��"(  ��:SI��+9D�8���(��C� R2`���d6D��R�*E�z]=��O_� �Ӂ!D� �D�S8vL.]��ά-�t�#� D�XpҌ],*j���䍞c,�ڥj"D��( � {�4��t >1���g=|O��y�GN�RB.�k� <������y�H1G�	�ĭ�Y�����3�y�c�*g�8�Q�� lѱԀ�7�y2�'n\���"-H�<	�3�ށ�yRÖ�2�6@�b%
�~U��ӨW��y�e��=ǚ�ȤƎ�p���#GI7�y��mÈTQS�L"o�v-���ژ��>9���yr�3��Q
Ή8w�|8t'ݹ�y�,ʎH�2�-��l�`/�$�y҆<>�p�c��� ZJ$�W�Z��y� �8|`)�f݄4�	��
��y2a�5�.4�W��}J�5:w%���y↟>f��A�fKs����֥���y��M��\;�mҭq6�;w�Ⱦ�y�21�ɳ	O���]C֪��y�*��Y���R�`o|t`�F�:�yB�	0�EY���ܦX�T	��y��R)WXQ9��^?+�Ĩ@$F�y"o�BԲ�9���<6\Q�R�J��yRJ���%J���)��`-�$�y"B
���1A�!�>u���	1���y��}��x�A͆0>��a{��V���'azBIۖW�(�C�%�~s�	(���y"�X#2+�xg��F�:@�'oS�y�	�8${�G '(D1`Fԅ�y
� ��E�q����1C�0h�8���"OTzv�T�O��-q�(иG�Z�"O\�� �oӄ��hRS�4EK�"O8�JџW�^�;�'�<M�@�"r�d1LO���s�8&珠R�6���"O0���e.�1�Sߣ"~�@�"O �#O�v�@i����)H�1E"O���Η2/�քJb�)0�M�w"OF���AHC����3Q@V�) "OD�#��)<�a�ML!.�q�"Or)�%o��ó+�\'�)�"O�$�C%Z�o',e��ɘ#QA0"O�H�����*�$K1(T
��R"O̐(&Q�#�吇f^����"O�h�/F�]�f�Ƈ;<Р"O����X�tr�0�fY�5��x�"O�$�ϴ�~���eR#S���d"Ob ���\}H�-N4T���"OZl�☥;�Hi�ĝYp��Cb"OHm�r��f��%��FRif$�a�"O�=�cʊ�_�,  ႎ*�.Y#�"Oֹ�"IM�<aR���D�1tBe� "Or�0E"�4r�9R��ݤN`��{b"Ot�q'瀫r�6�(ы���4�!�"O܁k���	�V�s
[�^�2L�"Oƍ�� KI����N�"ؐ�* "O���\�o p�I�m��>�)��"O�� ���Jq��QX% �b"O��K�`1w�|���	�u3�ݨ�"O-Xt�� ���h% eh�"OR��6o�;���ND8��"O�1�X�ln�k�.�%n�4�t"O2���]�r8���r�T�Xxa��"O�\�ѣZ� ���m\�0@:���"O[�F�~��m�V��x�:`�E"ON��Ɓ�׾x󀈞)~���{V"O��a!�(��di�e@F��)w"O(�B�ȝ�bI�U�E��&�zE�C"ORu��.$�}�d�N�y��H�"O��+V�R�65��jf��)��,�"O�E[�JF*j}�����*��1�2"O6�8B��c@� ��Z
SU|�BE"O��S�Ŗa&���p"�aXHh��"O��{Q� +�0�2`�"VO�XQT"OH䓣E�$�Tp�'�
9/P���"O�9#��".G�XI��X��	�e"O��)T+	�%v��笙�C��1"O�؀$I�G��ԐcI��ZJ����"Oj��w�^�z�*�v��$;˂d3r"O�H����I��-�s`�$� t��"O̻$�'u�H���{����t"O��)��1j���X��	 W�����"O�QA��9C� ���Q:�$T8&"O�Ȳ��J�v�1����!��!�"Ov)H7I �mA�yqR�ْJj\��"O��p��
�M ʄeM�zGx@@!"O�,���� �t5#@m�}�
es"O�qː��*f)�8��Δ`�@e+�"Op��d�(W+>�3�H�)��-�"O��W��5 bEy'��I0�3�"OhX�N�;Ƽ-&�bzy�"O��p�Ñ�:g���FP�-�
1�b"O
���!�jj	j����@�Xi�"O�q�7-4,z�����>\l��W"O� �1 Y3z���@A]yL�D��"OĤ"��A���͹�F�H�Ɲ�a"Op8 vi0N�B]��I�u��i�"O����ӭB�He�@C�4�ڔzt"O,�y%-R�|�Ј)q��9G�zL�"O��Bu�V�ZFx=����	+|��r"O���V��t���r!�?ꑐ�"O�4�p���\Y����	c�Tt��"O<���ٴ BT�����h�<)�K+T�jq�!*�;�A��Vg�<Q�`�;���R���]�"I��,UM�<�H4�t�3��8-f����F�<Y��'>�>$"��7oB��PBK�D�<��TȬ4��n�D����ECB�<q���;b8xzr@A�:>DX�4�M~�<�1Ƒ=.(4����J��l�2$�w�<!��^8A*C��7�J�#�'Ws�<�/\��!�op",�e�J�<��LB:8�(u�����O�5��NH�<�P萀#ߎ���Q�p��lX&�E�<	�a�w���`!�ԓ	�zc)�B�<AH#Z�p�P@��>>�Hd��{�<��K(B��H���:^ڱ�B}�<�kV6�X�)S)��3RC�u�<��)��_jNĠv�'2��A{�g�<�
{b>L3L�>��� ea�<�4KآX��Pw���w���
���h�<��'E�"�URF�� ����6D��;��W3D��r�[Z��a��0D�$��+[��آ�n�)5�ı���2D��xl5���BJ\)80��"�"D����!د IlL�҃,X��w�5D�(s&�ݚ_�RvCG�����3D����#��9��p9� /H_�� ��$D��Tl͙,�(�&	��j��%� D��8��0���:��IB�ߑG�B�I�=��Y�G0dT�|����3��C�	�jbY�>-z�b`�p6̩1�'rX�I�!�]�PR˒�n��T�	�'����C��m*�� aO�_��x9�'�|x@���.��%0�,T=:�
�'f�pC���xV�[��-JF�|�
�'ozi��CO�]��; ��E��e��'MDh��I��w�"�AwD�P�Hɳ�'�V�0����P'��x��߫@��}��'-�q��B5�᧭3���'C�z�aٴ^f�ٰ+�2�5 �'.0�joX
T$��@�zB���'N��F$��6����A�f�Jh��'��㦂�,n�ȋ".ıW�,%��'(&8AV�Q*Ys4MA!/�Y��-`�'���@ �ܪ8´8!AE4Xg�5��'�֐CV(�?_���#�%��h	�'H�s�D�m`!#���)�Z���'�b�#���$�`���ó%d�0�	�'���t�8byQ.4�հ�

�yb��=-�2�zWk԰�#T���y�� R*\T9/[� �b5�b"�2�yҨ�9wd�R�\'��Á�]�y�C�4**�Z�Dث0f<rr��yr��=�r(�%��2w_rh!1�yb$�k
�1���{����h �y�e���D��g��rᢐp7�]��yb�T.=��{B߫k����Ǧ��y
� U�J"3�x9j�
C't�$̲5"O�0���ݥa0������o�\�`�"O܈�&��s��8�pi�mȬ�R"O<uб`�F����U�:�����"O̩ٶf)K�����hĶL��5 6"O��
�"՗f�y��hBA��'"O��'���x�(�ț&X��"ODٻkP�2\L0�U�RD1��"O�)S�cY�?Z�{B��J_�Su"O���r���l�
#�ıiKԅ�"O����� ;ӊ�:ZG"OĸQ&O�D��	ӸrV��"O"p2�H�:�z��%!ǒSE`���"O�)�N�#gX��Æ\�=ȸI
�"O��dJ�-KT�z�ц}�$@�T"O8Ժ��\#fl��jRJ�`�d�� "O��vC�*�(�#	!&���1�"O�(siS���TGW/=�LLq "OPPK���*�d � %�X9��"O��Ǝ��2d�U2R�?��l0w"O���!�QR����40��%p�"O2�:��U0���n��	j	�"O��+'��8}�$ 6E���C5"O�mK�K�r��h#̎�K���ہ"Ob��d��1kdV�a�>�lY�"O(�A�)Y�
Xh�-M�O�l�ä"OB\�� 2$��lj���.�X��a"OF	J�pI��Xp(O�W2A� "O��ג�Dq���eE�,:�"O.�be�T�U�e1��)Պ��"OmQ�N�5���9ŎC��P��"O|����݃>!�!�P��L�R�Y�"O�q��圖;`�(���#V���s"O���֬G/"��a�`0��z�"O����A�4��
Ԕ`ڵ�T"O 5��)I1����َ~g��9�"O���$˺/a�R�N�r���w"Or���B� ��5�m�(^�2�Z#"OΑ{wK�i��	Ywm̝;�,a��"O�A��ޙz@���~|Qc"O��Bb�� e횔x����K�Q#"O�|p�ӴV	�)$뜚@�n=�"On)Ĥ��d���*Q!#ޘ���"Ob5��ٱ&�,���cߐg��s'"O�<�ЧTaԦ�ЖCY3��$p�"O�� �A�0th�F!�8lǖi��"Ot)`�e�|#���A��
��"O8q��)(�")z�*�c���"OB���ܔ�6a��#�|J�"O (�&%F���${���'�
U#�"O�P��+�����E�4)�"O�����!�j����5#p����"O�mC�(B�<_ ~6���"O�ՁF�ߢr6ȹ�DB[�&�~}�"O0�J4e�*j�J�h6��4���g"O�"��I/肙��@�+-~i "O�!�g�[�|gZ���n߈
"���u"Ó'%Y�&{4y!��ۿ^���2"ONXy�#��<lг'���̰;�"On�s��#4kb�:e��R������':�'ﾠ�$?%p�q��R7�P��'��)$�τ�#�E+!F ���'j�X3*[�]Ƽ�Z�f�b� ��'�F�+g�<:�y3��M� P��� H�*��:�M0���7�|�ce"O�T�Ve�JU� �2AϜ��A��#4�|"��'l����i�7Dq���*D�,��I������p&�17��ҟ,
�F|�P�$�R�W*p��ݙVPt#=��T>5�EJ��u	�z0n$��l J#D�@�t�$H�r �H�z��F D�����;�6��U���<R��?D��k�B^-
F�	�fgQ���'"D�!�h�((��xsΚ�O<�a�)>D�DbH�>\!X�[��>i�b���:D��hc���#7��Q�FA�L��-D��:2iٺI�~4jD,��D-6D�p#�!�"K]l����iD�s�5ғ�p<)��ȉM#D�ua�7�i����f�<W�X�o�� Rp���r�2 C_�<�@�-�P�X"Cg��8�O�s�<at�B�L8���@9�`E0��\x�	c8�$��/G�y:���=�L�� �O��	�i��$ 2n8	�%:��05���'Qa}�
���Q)��@�A*��l���?!�'d������6k�9K��F6!�����'h��Պ؃& ̵C@��I��R�i�F����Y��,\M�i�傍c��B�	�yc�\⁄	#42�*��0��`���<O��:�*�h����
%��C�"O|�4A!k@"i0v>�8�"Ob�ceY�@��CO�:��G�'�	�$srh�4�چi����S�+B�I�] ��ۀɃ�Z�Kc�]�|��C�	��Q��f�'p����������3z�nu��$�0W��ʷo'	>��ȓ��4K��L�u����FUV0��8y�ma�)�i����ah��w�����hukK.1���2F~X����	K}���M��$��mP(0\e[7gϷ�y�j��K� Yӗ#D;�(Y�	���ybD���|Pee�$y=�e���B��y"�L�H�;T��tҚ��C\��y�� 9|<p9�b�> U|}X@M�y�7��z��OC$ `H��]�y�͒��\uZ��	o�0�����yb	Z%)� 5�"e�*�Q�Q�7�y�d׫"%h�+�Z|əj���y���hԊ6"@�tFB 8P�ۦ�y��%��Cc��7 Q��&"֞��'"�{2c9b���H'˜;|e�Qv���y�fC<3x���J�tu�P���y����%�8� �	��=A�yr
ϾV#e3F���Tǂ�1�kC��y�JJT�%ʗ�٦R����iҬ��'x�{�쓊��8��ΐ0NK�������xR�'�� G�M(( �<��_m.����'U��B�)
`�jR`��16(����0>IJ>�����$<�+B�J�X@6q�r�\\�<����^�f�KkY7F�:��p�q��'��#���>#m<�(%�X�m���j%2D�KU�I҆����Gڼq!c0D��k��++m�pe͘2��|���.D�\�O����=���==:I�n-D�@r��U�'�j��e+ײ#��C�*D�pH�%O���(gF��f}�k��(D�|���Ж&\�pA��>�G'D����H���!s�Ԥb�D1g,7D�� � !A
�"�h�^�Jc�9�"O�x8��N�y�]��GN5XIH�OH��U2�+��ʞ6sN�[��R�D͉'�|�̑?;k���C����EӈԨ�yR��7g�8ȹ�K���)�R�O��y�J/\f���Ry��D�4����y�Ϙ�
��ݘoN B9�y"�%-U�}�s��u|�(A�!I��y����8�.D��fȚ��t�N��p=��}����V@���N6�2ik ��3%J6�=E���v ����T=�r�y�K��U����=9������"AƩad�|�qH����?��'U��27��*њ��&�A`�6P��$1��t�	�0.����
�l����h.M�B�I-`ʀ����Yr��?L����F{J?�0Å_*xu�aX�7f�u #�=D�����I�Mp�la� :~��-#��u�'��#}�'̾Uk�!�%U���T�����!��'������5/�|�h�-lĄ�{F��OPC�	(��(�Bk_��Bز�#�d�xC�>g���XDo�F�i2�Q0!��?q��鉢N>T�C�V��ņB�&e!�$C�W�rd�u��-�Y�Ph�M�$��(O�>�1�ɞc�(�d�ڠ'V�P � ;D�TPt�X<6{�'�Y#�<����&}�Y�؆�I�Y&,�a���x� ��R�,B��>�}Rf猵3�����b/N�E}��Ӽk0(�%+���M�P>��$1��̾w�йy�9b�fq�C�++��$1�OdH)���qIm*V/S�ms�1��'�1O���$��$C�\��م$�I��|R�'fr	#BΖ6�2�r FC}�H�(�}b3��?aBP�হ�FE4( "����f�1� @ D���"LQ�R�Fh�e�M�w!r�jD��=�M��{��i.��b��O��}*�>R� �*�n؃Z��Tz�' ��V�'Y�<9���Z<�r�'�ў�}�r�Y�*ڴq����MH��b�<�fe
=���2��M(w�^92��Wu�<���C(xS����!T�`����j�l�<�CCW6N_T:��䑶ET�<�,E��?0 0ʰn�� ����AON0$���(=����"��*�ȑ��%;��C��+�z}�!F^<2u�ay�K 12�C�I7B]n���׿K�:��&з#M�C�	�<���R
ǯ9�@LI0�έ^jvC�	�s��� B�ԭi�T��.n �'������R�6x\�����O�p���!�R�<�`�O� �|u@b�~Ǩx
p�I�IN?Y�{��$��@L�x�Bb�9�>�k�g��l�!�!yԶ=Sץ�j���8��ק"��M���D)�	1���7(%�BP����#^��C�Iܟ�z�'E��	�����:D��#R�W� F�U�y�5!��.��%�S�ݦ�B�D	�@-h��m����!�9D����1���5�C�N�J�9�6�d�ݟ`�'��3d/P��vFUk�,z����}hC�	g�t8�b�����v�NC[B�'0ў�?�*���;�:|���	W����'�O8�'�z$��,����{���x7\���'��E�e��L��3�/B4^p�'�iX��B�4*Dp��3�Rda�O�� ����9I�`��X�$�F��]�0Γ\��In>e��끺]e�Qw펯Je��+ū>D�$��h\�
���R��B|�A9�H}�l���y��F{
� ���ܼ[�fQ���f�x�+�"Om�D,�;Rb�-�q�Zo�~��&m:4��{E�]�g`Ҹ�V�\7d�P��'%><Oz��?��ρ"q�%����".��U |�<QR�͝v��pi�2Q`�X���R�<�阫��*4C�/�}�IY�<q�gʺly�ш��B�!X�`�A�
U�<L�>yA���2WԤ5P��f�<1�fS/`���N��{��M�cz�<ٶ!������=p�l0ڣ r�<�(�����G.8#�I�aDj�<����R�1�k@,�t�AG�h�<a���=~���K*b�F�A%f�y�<�SD���i3�� ���Rc�v�<����7�&
�GR�nAP�Xs�Fu�<�o�(<�VHГ��6�H@�6��{�<!T�� ��R�@Ҍab ���|�<����-#䢭�-Q-3�6��	v�<����p�$�Ɇ*�"Y����K�<)���>fu��"�
.Q�9Bn�n�<!T�G''����Ҋ
Q�(ę&�Jk�<���S9?[��
���7zD�'�B�<!t��tZ�@���.U�%
���t�<����d�Μj�f\�R>V83���f�<c�~��Y���7bI��Z`K�^�<�l�0�3�(ܳ!#Z��U/[t�<�&#G>d/�Ak �������H�D�<9���(�Q6�K�X��P"��w�<����%c~PR���Ha[t��M�<y�/��w�l]��MI�kC�H��	`�<�vi@�9��Z�i]:z��m��d�<��i�q���"G�ϸ��\���Hv�<)W��%ݸ4� �0�R(q��g�<D��+t;���a���	��$1S�{�<	��-o�y�I�3�^͸fM�s�<!f���.dV�;��Y�r�*�Hf�j�<� �?w,�0��3L��y p�y�<�ÅRL �j�&�08x�b�O�<i5��)��E[��A�H[X�4��E�<Q�{~:H����"�&���\B�<I�G��
��w+�8��A�y�<�)�6b�y��C�q�p8�B��B�<If G��� Iȉ�I�jIR��Gx�<�n0�Zm�Gό?�X�!d�y�<Y�LʛfK��@R�S�)$h� �w�<u+�U��h�wB��xD�Qd�Hw�<��#�-69(E�qA
=��(h�J�<1PF�uؼ����c�:|�"�A�<)��H�b� /��
Fx�y�D�<�L̳q��9�t�F=���QW��Z�<�1k��bJ�\3�`�	\ԑ��Dh�<�Ek��h���(�ּ(�e��+�m�<ٱ�V�QM6� GſMV���%�m�<A��C�rF��(i�Hh2y��Vk�<)b����l
��hi{�<1���@�!c'��&��
#s�<I�R�u��8�">}��,����n�<�p��BVEZT��~d�ѧ`P�<)t�Naj���L�7uxy˦eu�<�e���)3BS�D�nӃ�s�<i���59lXh�*҄=�eH�mXt�<�g��x�
�E�z�N!�$Wq�<�7�	*s(���h�\бJ�<�U�?t� �C�pR:}t+Z@�<� ^`�b]<l�bP�s�6P;c"O��j�&٦JQ&|����.l舡��"ORe1q�I�'����JϥQ��ū�"OP�cd��F�A��D'=�&�@�"O�H�`)R5nr8$�(Ş{Ķ4"p"O�t�\�ޞe�Ƨ�l��Z`"O�,�q�Z3��1C���F��ݺc"Ol51T!��w��\`4�
�j�l���"O8�2��s>�1ӓ��&E�F���"Op�`-E�z P,Y�L?_I�"O���؎0���b�3~�����"OZ�s�,��&���j5~&8�`"O�Sv��J����3����<�"OV��1Ѥ�8p2���I���3�"O���Vۧ����uMV�H5:�{"O��
d���$ջ�X�7_�((0"On,rGn�&������3JL�-�B"O�}۔�N=&Ed�FnR�;9ԭ���'vv�K+�����Bʞ;�:Q�"�<@$��1'�?D�$�w����`v��T<QW�:ʓuW�1�'���H��Y#�bH.<a��S �¡g�Ig"ODE��!T�oULŸ`��9I����dԤ	L��6e���)��<A�o�%9�(��ǋ�wz���N�<��)�3iU��s���x��C���<���<�t�Ȑ�7\O x07l��#�>���EQ-v���'�`���H6�FJ�IC��07i�NTH3 R��y�O�C�A�j�"O��D�a���O8��Tcʜ �@���N9YڦURbj�p�v��4kMt�!�D�3'��AkQBO��I�ΈB�@(KB	�/�pI�"~�dw4�9�i�<�R�`��.$F���$�	"kP�h�5�M	����Γ!�
J FZ!ݐ���Ƒ ����jH�d�h3#Aa|2��z��8� g4p����:lU�L�����F!��'���O�F����fҪa-:�ʍ�Ө^��1!�/�'�LLr�_� Yvd�G�(e�P�ȓA�����+F�Jڼ�0�"G�l���n�75{|͸E��sӨ�`�66�����S�Uf^<�0"Oz5�����"�Q��8,=��"O���td�Yb�9��`ӡ2f��"Oh9���Eq�b��J�e�"Ol�d/���`Y:O�HQH@�O���f������h�� ���ݦB��u���3zbt�"Ox�원Q�P�C��ON ���T�@!biO�|�61	ϓ,��Ȳ'&<t+��G?�t��I�7�X����Hg
������X�RU����9N�]���@jH<IC��8�1�l��yi0�P���P�K4� �FZ{�R�e9��0���1�-C�Dc�ף���PB䉻Wڰ���ER3Jޮ�B�CJ3M@�c�˹P<�DJ)E?�D$�g}B�G�1����v�W7@a��9�yr�	X���P%��	kqlP�M+1k��,�8��"�"d*��	�lh�#��Ŏ�H�� %E����	�"!��A@H�bd�!���=&���r���3nw����)u���s���.6a~⯟3;�: �  �(ĕYui���'�̼���ֽ{���u���LT�p.L*��iW$F�rF
��,K��놨�F�!��nr�T:g(��:䅏�t4<�0���4T�3�Z�@Y��aG�AB�>t���;Y(�`g���e0\����M�T���&ʑ��R�<�,�@�W�����"�)*�8���N�"
je��ϭ%�b�I=]�X��ٖ 2�w�%*���D���5aSn����Gl��`�����ɦ>�B,R��X&�Xv	I�>�d��I6R������ �4ə2��$�&b�́rD܉ �0TS)�>�z� �R�/I��X��������n ~� �(�2S���"O̴;�e�2H.D����%f͎	 w&L�QN�4[RA2LYueƼ�~2 �ؼc�ˊ/^H؉���	 �\[�m�<��f �L�%�3z�h��0�׭EE�;��
Zn�ǈ9	[l�
Ԥ���HO� �ѓd�܎D4�	Ң��?e�jE���'� e��%��L�4�1e���@v��ȕ�.]� ��Q��x'
�R�R��2�OzT��%)�� �ɐ�j�$D������E.ջC�,-&<UyVF (O�vEk4Q>=��*@�g�䔀��S�:��T�P"+D���օ��p̐x����CƜAG��n[F j��I<�q"�!L�u���|Jghi���3��4�N$
�3:�����:D�@Y��}�v�@�KY'���kv�nӸLB�O�Df;��~�,��D�R��Q8SMI3K̦}	�MC�9]a{r�4.�A�'
�?�Pq����[��u[BN�2Qp�CpȗL�����"v ��"-��aZb�9(�ON�2��5O�`ңMXV�Ӥ�~B&H\1�zT����&��Ȋ�h�L�<)��U�h�"�	-u�����U�Bo<E+!�I'R)����:nZ�D��F�"�������$ď��f�b�� D�4;ċ� ]��5�EX9%�2�;�(��@�l�%�[[a��C�l��0���g�'x^�����d��[��<4���
�4����U	�;C�:>T��e�!z�J�θF:���c�'��	�D��TP��Ie�]�	�3��P@��-?�ʓ=t�\O��
�b�xE����"OHI�6f�$LV)Kt"�e�V�:��x�H�7U�$�J��i�O��x`�cŕv���PΖ<��+�'�����ϰ`(�EK� ]��bVLO3�K�d)��x�cG'84��
�xmbt���M���>��ͨR=t�PR�])}(l�gjY�C\<��)�"CSȽ�w�C7z��}�I�?�t;2k�
r⭈
�HOV��ք�S���'4d�1�.��T�4� M�"��̖�@/�,@"OH�xEU8,����ɕl�����VQ\��­� +��L�n�?h!Q?��ܧ3��D��ɔ�I����d�\�LI!�H���tA��	xP��� �!��4[�"H��A&\�"#�?�=���Z��=G���#�6�CPb
N�'$���E�L�䒇qR|��	K�˔I"A�B_���@7�گ8q�X�'��[$�D�����ċ4�ѤNX<G7@dz�,�)3}�p����9��q��3<z0���e�[":���"O�1�F�X۴Q���V/��3�șjbj���|^���uW�W[ܺM�W���
KʦxK�F�l�8��H���
��G�ǃ9
R6퐷j�v,�`d��6���S�`\  ��$� Sx��O���0=��fC9J��|�@��"� h� ��k�l
��Lq��j�}(� ��7ȥ� �gφ���fZ�A�Na�o3D�ȹ3
[�c�Ԡ�DE66jd�+"�8���[V�M;��d8;rLu�W�=�������-y'xy��Ѩ=F����&�q�<��A�LRI�Wo�9�$�����$�~��m�C�>b�(��c�`2��W�8��3'�!p&X�ө5|O�=!�'<�Vq"�4o�����Zm0z���
����f1<����
)ʁ��A,,5�O�B�C�+=�R@R���"}�b(O�=5��;6n���: ��m�g�<�e"M;FZ�������H�k^$ڠK�%�?٠oO6��Y�|�<I�%�1~���3A�)�D��c�In���Z���6�6��&�O	0}��qQF�=��$SC��oc����X������dPm�����8���9��r\�E�5XlL�N5{�#ɩk���J7$�;a�l$[�x�.�6v��݄�	.'b��FK�yr�t�$�Z��H�,���I)h�	�`�`y$_>1��W�<jP�1	rޱ�Q#��Ա;�)�cH<١ �#1Y�kp�N�K;P|إ�S�L����c�ZV*�с��2^�CP��I<D�i�=�6
���m"�O�0�d��'?�O�)і���L�2y���	"wT%sS�4.�I���S����y��T�vt>�`�B|�l���"u^=Kg�>)��D��ݹ��D�H)J��L�t�'�=jק���*���3ԚP���J~�Pb2!b	���f�G�zƸ|�W:Ot6��h|p�ǓkT�vM�E��M9��\���'�)�G\�)t��I��m#(�~Q�IW�B�^�1����p�eE��Zd��
²b�t`�'$��𰭂o�&�s��зX�tmrT2O.��V�>!!y����'F&���p-�j�,�s���6�y�w�l�[��3'70$���(�'7̥�"��9���%&��.�2�SA*��*��Ӱ��*\j�E�b�:�8��SC/�Q�U����]�F�6hb�`��I�D-H�Y,#P�� bwZ��@G+D��"5O�IG�~�JǓT =���Ӽ1�1��A<j�d�D}RE��z�6�+、^?A��(�� F�Dn�5@���ǌU�pP�"3"~H<I�.J6C8�X���(^�mrBfOX}�aųv�L���\�@��&����~�*0��#<�@Y[�o��a�l�jU"Oz5��#�)$4ވI�G�%�^��|��ǋ$�Z����(T�r$��\$r�k燐�72�l�	�':�x�ӭ��"a6���Ǵ'>��	�'�V���P�t��ҦL�5��	�'��ap���x{X\������'�dy�C�^-l�)õ�������'�Azv��&�8���ۮy"H��
�'r�x5��#4�uH��E�\�	�'�$D��� u��#�a��0u�u 	�'�� ृ)j����H�>}+� D��
&��X�n���`W�p��+��>D�x��Mƫ~լ�a�o��إ�L:D��ɀ��6A(�@%Eݶ����;D�D���A
_��Eݟ,_�����:D�x���Q1/�i��h��
3��8D�ܲW�˳fج�� W9Q291�6D��f�L��!Z�,���.��(D��f�T4	J�P0r�� BhZ8��� D� ѧd@����?4��{�%>D�`���1-���Cg'�(b�X�[�!�DW*.��`�$NK�f!ѧ��!�d�� ��H�U��5�v�k�F�8�!��tC��v.k��ez5옸�!�D�?,����J�8f3u눴R�!��{���b�m��j��!��C9�!�_���ZǇ��v�v� "%U�c�!�$L�J��H��^<vh’��_�<u!�+LH�P�eҏVkT�Zv����!�Dkql�@���͔�hG�4}X!��C�%=�@Kw$�9'�t�z�N75�!��4	����`�&$i0n���!�J�2�x�z��M�}�������!�DU:J��EI�7��'Ά��!�$52�ޕ���	,��UKڍW�!�$��&cr���bg�@�j[�z�!��(z�րpg%
�BBv����@&�!�$��HA@�y�&/�y������!���f��\�G���#�6�#��\�@!�d��
�y���R#�"�2f�"�!�Ч~Y���$������68�!�Ъ!���4�[�k�
$���/�!򤘍��=#�:U`�G��P�!� �U�����	\����M�p!�d	/[�:���d��=4T;A�[-j!���2���zf���6����.j!�:Jo�@�5i�24
�)�"��!�$*��J0�.�"R���!���4!����Fp�8h(�E�!�]�x�˄^�2ؾp�ů6�!�W�4aQi��(���T�G�!�\ Dh�sfX"W�")�մP��"O�<���
�0D.� ��#T��9'"O��(G����!�'�28�zd��"O*��q(B�w"��d�9e-S "O*�y�A��`�^Up2B�e���"O��Ç B� ���s� �1"O�t��N7G	��@�.&#��Ȩ!"O ]Aa�%��!�O�����"Ol�D�:�p�.�*'��ؐ"O>�@�>_g(Mb�F˃-v6M�"OF4�#I7,u���&�,Qh��*p"O� �a�#-�RfA�Ǎ�&f̱�"O��h���!��u���OnXxy"O�0ƃ��0!��䔳[Y`�P$"O��蠥Y�CnB	���B�Y�U"O橸0�F�M�#� ,1̈�S"O�y����u��x���ؑu�D�"OXTj��,"�ʷ��5V�b)�A"O^��c�J+G�dq�E�?V���P�"ORy��	�vB��{�A�&���#"Od�I�Cُ-O�˓��jΠ)��"O��jƄ��-}��F�	>P����"O��Ks�K.��W ���%I?0�!�l>�(�@ �H�(c��N7p�!�F&|�2��s�F٘��G�!�Ν��x���>{�Ih��J�!�$9����7 B���Qψ�B�!�Մ[����f�T��r�ג>�!�d�2|�5G�b��,�@�S�	�!���=�<pa�b&_����"֗TC!�
;�,g�I�/�d���J2!��Rv,�����Sqn%�Y"O��+��E�����F�o�)��'��B�c������!G} 	0M����b+D�Hq$"F�{�=qC@ә6���aG'ʓt|\Yt��
�H��̫$�
e_Zz��c���0d"O��E(G�> ��[�&
�&� 4X��J�]�|�c�8��)��<�3"�HY!�</z�EK���V�<)� ��En8j���%����@�E�<y$��S��kҮ.\O����`<`*ڑ�b͊�z�P!��'T�ȓw :���b�$�,\��8"��^x�i� ���yr�uHHd�2� �,Ȉ��8�O�l;�f�8 ���؊�J�-:p;V���;5M(U!�d�� 8D��f.\,p��*�)ژ93B,3"Å�l���J�"~Γw����EYm�z\s��6J�J�ȓ{�0�a*$���)3K\��͓Z��R� �	)����dÖE��#��=^ (�c&$ka|Ra^2Z�V<i�!�"g ��%G8�FY�TAF�W儬�
�'�X	�*̅s�fT�#����m��^�< �L)�
,ҧ+��$�2A1 !3�+��0,�ȓ\��l %�ԧ]5��	E�0�r�lZ��@����s�4��&B Ddp��h������"OL�)�j��ME` �'���ر�`"O`x��<�$�V��Y�>�R�"O�0�+!Pb��0L�� ���(�"O&=K%��5Jk�Y��� 	���Yu�O�YJ�������h��!%���R"�lB��J�}�<13��	[���y'`G�{�dy"s Vu~��.�~��T�'<��P�rw0L��˜�8�fk�8�lS��ک=2�j§A=xazL��πo��p��#$����'��\Ѹ_����e^�\ўx郭�"?���Q���tl�Q���W*���cϿv!���Z%"�{S���5��qZs�.�r�B�2���o�g��S�/��ㆍ�B�P���S�/�<�ȓ.{���qoU/pGȁ#�h��<��'��q�n�\2<��	3" � ٖk�1c��K�Se����7Po����dK�w�ŀ	c��VDBR�$�[�D�;{e\���k�4� Ƀ
-�IBY�Oў4���?G<XҀ�˪G@�X.�,<��ۢ�<H���4���"O�̀dC���,B��9X�p��'@2����#w�4ݩ`U
D۠�D�d�,�]@��=��kq喏l�!��5`,,�ԯѶE�t�[cAX�HtC�ABҦ1����|o([��"FxR��"*:�e����Y�4@�.�p?��ԁ
��PZe�7o��M*r�S0إ��R$V��A������>�M�|�0��S.<6�iWgx�8���R�0"�Aw]�� �\!�?'���L�9� ���"O0�y���,&��赫B8�4 ���'^�rB݁^� ���1Z:�E���T� �Ҭ�!��I6��q%P�N!�@�p@�`�B��>^���X5��Ig��V.|���c�+��S^?#=ѕl�>g�i2�"�
�|`Ɂm�^8������7f|x1K�=u�}K /V�d�C���@Q��c�(��f���I�hp��T ��E�)H�L���<�t�I�mz�<�`P��Q�Ci^���]�C�2DQ�[hQ2,��yn�0.l��t�F�[�����$h�2�@B��M�d@��	���D����'� �W.I.xZ&]1���KRP���'zT�9`�ʕf�j� ��K�O~�m��'T�(S�*QZ�u���#ap�z�YN�|BsDοk�p��D��:��U�'�m��d �����B=&�J�'?$8�>0S�|8R�NG*v4K��$G�G70X���?1R�t(r�D�)
�%����c�^$�t�fG�/w!�D�)8����I���;��"t�����,���؁k�0q�1"��O�Mۑ)Ԏ`��AǗ�hd��"OLE�,h��X9t�ؖM���U$�5�"����Aeє蟮[B�3�v6>a�7*�/.@���XJt��	~N|pw�''����Ł5� ��(�M�\�CҬ�2/VH��(%4��暑0�t��#�ΖxE>���I�!f��:�G/��		D�Hc�"�n��-qY�C�)dI"#q��8�q�1�OtII�c� i:T#��I�E9���X;K'
�@E�W�!�$�Q��I��FP�5-�I5��+J�
�)��>}���R�jc?O��Q�Y+4		�������i��'���y�_tĎ�����5c��X�.C2@�rQ��(I��}�?�O�8p A��:�|q��M!��<y��Z,���Q�4X��C�``�S�?��P�"�#?i���q�J�m��B䉇Hj������u��(�L�� _Hx���<0%xG�� Ȟ�)Х$��h@d�@%N�nPv���M�F`!Bh7D���f	]+db�`r'@�u�p=��DRn����H����n�.'��@�g�'Ķ�����x��1k"j�]�092��$#2Ʋ��H�$ŋ%Aj�qA#�	,,H�Ȳ4��y0�
�c
�J�!��1w˖�H�/�P��"�Tv�S��I�v���5�TP�X���c>�]�7��1�wǂf��@bj��V�C��r|Xec�C��"�B�w��0�GU�"�&�(0Ό����ZmK��
��b���T��<l��@s%č���@b)|O��!!,���4�T��6��09���c/�U�Ɓ��p��1�$Nx���D8h^����'B�2{�%���׽	*�O�삗��vڲ��)O�AӃ�\�I���W��"�H��yF�ܫ�1�y���z�*��vGV��|�qҊ
*�h��lY���$��bK%x�.��|��w�1Yc��T$���y	�'dE�!�uӺ��������E�1)�Z�([(�'0��sr�[t�=�. �#ش(��aa��A�}����T�\���[�?̛�oX��Uhc�֦U��M��iƭ�y"&ܭ7̝��eX>H�n �I��}���" �	kʘ����y�O��uB���+G���M1K��PI�'���
g�\�T���OGur�P�/�*Ru|��%�'���Y���Ϙ's.�)���e���P�l�\���\q$��ė(5.�(qL�.z���+5��CNr��r���P��g0�2Bb�#Ů��� νE5�%FrH���`<���WC�S}�X�׈�5T��ذ�]�p�TO�`;�!�;��<Ya@�-(�Y��̭<�
!�q�ZyB�7���{�lFi?�%!
���'S�ظp@֌W"FɑB�T>;L����V3:��p�',X��f и�\�r��&Y�D��e��ːhU�t�RM��-��-\�����X�b�k�d?ͻ"1���t,@��N�YFI�1N�fU��� 6��ɅFS8^����VՙQ�Ҽ`�*�Zd ��E��l�@�Ո
5��̓\��DH��R���'�v�Ku�� d@Y�&[�y�l�)��dլ!�n�������?��g@�X�FA���Z�m� Ad�Ō(�Ak�N6��牐F�L��2�5��x�j��`Bq�i�ĝ�����d�$/�L(�"�?	0�X�V��h���`>)B�CR)��MQA*�g�,�C��r���������4�2e�4�ݒ?N�UIb�Av���&KT��#�$� a@�K7�*U��E��>N�]i2;O��R7bl���Va8hg��#\�����1�� Nt��������� 
D���U�ķnh��q,�=j�0�/ɭY��ԟ|�I0�a��?�\i�����18nD&Ax�~�ɐ��4����}dc�����0lܘb8Γ&p���C�3���D�c�|+�Ǔ%.(#���2N3Q��+61a7r()A�O�y��0AS����Lޜ.%B��X9��5��($�X�W�8{�Er��ӌZ�.���>�s�҂�n�b-O(h02'�9��O�S��/H����xA���	�'�֘��I�l� �
t��~��YQL>T����F*�dꢁ�>5о�2��H�@i!�^![�ya�!�e˦InM�n�!��*=��e[�N�F4��wbM!�Q�Z����2��G�]��o�5B!�	V�rQ���*Vo�x����L!��$����H�Y���鷯	�o=!�	1+� ���!�S�&?�!�䍙q�2����<M���qa��!�̥Ş%9� ��+4���3^�!�$X�b"v���/=4 <�T	�~�!��Ęk%)������	N��!���Z��J;T�R� !��<,P}a���jȔ
#��0V�!�d�8sX�eyf�ީj���0D �)�!�dY�R�p�8.h첨�%��C�!�$S�'�L𢍝7��]���ɸZ�!���R����L�BA`m�?5�!��T%Zl ���3$c���ǆ=�!�$O�=H�䫐$�!��835F�-�!��ђd��͂��C�UU"0���Ac]!��Ћ^��14�Og4fe;C�rO!�$����)��/UY��h��Pyb�˧(��VGG�[��+�ت�yb'�)^�.�#c�{�����y��N�0�z�"��pK.IJ�bG��y�D�ZjTkF
X�c��e��yaPH��#ϑ�!���C��с�yr�P9j����o���i����y���	z.!�H!\PѲ�?�yR�D�4g@�"
��$hN����֤�y��$6�<;'c�R0�'O�
�y2mQ!C4ɒ�'[&Gf@���T�y�咺K�2As%j��?��q���*�y��Y7fD�$y�mڟ>||;E���yB(�\��I2��< $0���y��P����ϊU��y��'�?�y��A ?�@�p���HON��6���y�A�bDa��Y�2�%+����y��	��pC=�ɹ��Q�y��Qu1N���_�D݆Q�����yB�E
 ���<mJu���C*�yҊ�$d�l�����/,���UF��y���-rF���ɞ �P�:4��=�y2�@�@Z�-G��Z�����y"B qw
����I��	�!�'��	�~���O���Ƨ�yr"×GT	H�%E�z������=�?!ad� d_P0P�G�����>�ꖅ~���b�t�RY$L_�[t�t����)��p>U�n���4�*����W��Z��1�j�<�&+���i+ba���I|z�M���)Ђ@P�&o�a�7��47�VL� o߂-	Qc�&\�|�ZH��S�"�`J�ΉR�>y3F�1c�F�20BO&dp� ��ӷS`F;�I$���(seFlp@���}M���D/v�<�:GF��U�����ᦑ�Վ�G>y�df�#����ϖ!"��T,�'Jg��9���������8��!��=<B4� � Ǩjo��4�(h���3d��
r���f�H��f?����� �<z�u�PL� z����?�̫7!�
�F�X�ר�Ң|��O(q�g�N�^4�����t�^�ڦ�R|�� ��aþ_�B�E-�O�O��r#LC��j���/nax��3�Y�7�60Ƞh�,8����0|� ��1`�"6t��pg�'u՚���e����(rcv�yZG�I~]a�T΂VS�m�U%J�8���jCV�.�h%Ŝ�XT�0��A_�9�4@iU�"�'�u�&g��UCq��*��͉��a��hz�	�V�ԡ���8��������N=!~��&��)`l��iժ��2���jS��
�OT���>�r�i_k�8�AW	�?E�f�ϩ�y�
Ju7�K�@��-�dD�p�œ�y��N	�U�� �BIY��*�'��q0�`�A���(E���sO"d�'�hlåF84"���t�2z
.8��'p��Y�� 9�^���ʑI�^���'ص��˝-J6�]��Ԫ<���
�'ɂI�Ѻ���1��H�'�����J���OI�8C0���'[:�ڃhM1��0>l�q��'7�؂!�	�p��ã�$�ĕz�'�ΝZ2��}��s�޴~O,���'��B�GN	71�4ifʬv4j���'=4�����8��jb9p���`�'�Z�#O�7s	���rK�b�@ը�'Z�tӃ�;�
�H�+fN���'d�)�WJ�:v�s�Ì�*����'nxa�/��yg�預��#j�p��'Y(��C�,w8≳�ΝJ�����'���e��:|ntA�c�z<<i��'�xT3��I�t��;)M5�l�B������Z�J�ChJ�O�. iQ"O�|X�"���~]��:N��ɰ"O�e�F�/�]�SFR{��B�"Oʁ`@ǟ�Inmr�N^,S�`0�"O���NV<�D�m�D�lp��"O���!ͅ,�����٨��s�"O���C���`�3(���fx2"O�U`��/Qv<�Q��0n��:�"O$EyqC�L��r����쌻�"O�P0U�^�F{ޔh�S��A�E"O=S���|���0��y��U��"O2Qb O
�
�� �R �B��w"O���EI;U�Zak���2~Q(TCu"O�W-ݠ2ʎ<�ѩ�	5�z�Q�"OvU�#�� J��]�gcT�m��<��"OR�) �д�� ʄ�E���!�"O���G�����y���:��-7"O0�+R�C;RT�U�M��J��@"O���i"D��s��X��y*�"O� B� !���X���.4��*�"On���߄1�z��B�P�7"�	�"O�%��"<NXf�""��;�1s"O�hhg�*�
a�Oz�.���"O���!�	i�*��T�߯>��Y"O[�w��N��<�flۑ%���;V"O&�d+��B���r�*=���;�!��@�4��Q'g�'�����z�!��	�	��H�G 6o|���NX��!�$�+O���H�)eTK&���!�C�F��D�F�qF@�Ӵ�U'>+!�.g�2x[#�߅1�1�#թ4�!�E�o]V�R���#\(◡�#w!�䑆I<h�pG�&�<�z�P2�Pybký5�Jyc�
t������	��yr�5�
q{�䌏h�24�ek��y�/]�\��d��j+�	Bd�	?�yr�;�̸Pkτ^��rdd@��y��E�H(�sV� Z�8���ʖ�y�����s��9Sf��%bZ��y
� �a��]�/�<�S D$D���#6"OF�C$�=FL��uo\v�е�'"O.���퐱PgT�X���n&��z�"O�8
64R�L�#㠘�A!�}c�"O�i��.J��r r}J@r�"O��C��
�-���%PKL��"Of�BmD>X����CϘ�{+*��$"O�%��(��e�&����%�P��"Od����g��5�����2]*4"O0��Re�0e���+��C�7�P���*ON|(���*�l� �M�=���x�'���sJ�f)���a�m��'��t�r��#JY��F�WD&��
�'<�,�	פt��|��VJ� q�	�'UL����m^B�ٗe>�ձ	�'nd	Ić�?p�[r��6��1�'��( ��0>$pb�AR00K�	�'������Cfa8���0]�`��'� �ϵ ���	ԩY<Z���'H�wiB7&�p*5	��F�e��'����I��0&~�1�D�+2��K�'n�]���P�a��� C�+&�1��'�y�AbY�����E��tm�P��'�a�5'G;��@b���r0&щ�'-�yP�����J]$N�;�'�� )�H�/�%�d΋Wd���'���
�y9I����V�dxp�'[@����Ca���&O�N54���'�h�2#ʤGS��Gh�$M�
�'���h3�\�n�&�8Ů��>n���'a"i���G*BL�������4�	J�')`�a4D2Z�X���~N��
�'�.(��Ud���r�#c��	�'np���ݓD4�8҇T�\:����'�(�2�ϧ?���bZ&d�����'y�Գp)��F��H���Z��1�'D���v��7Єy��bJ�	�'��}31�� Q<��ՠөm��-�	�'Gn٫�mі^W��xud�	gZ��;�'MA�Aތ0��P�����R0���
�'@*���Έ�H�x(R��%�x�
�'԰��2	B�����~�6(
�'�\:d��)d��X`�K���H�	�'��AK3u����M�)/��y��'�4M���~䁑F�۩y�z)x�'��E�c����@
��إi�2���'j�� ��	��,�F�#]B�Y{�'<�D��Nц'�h	
�	��=MJ]q�'lpqK6�_�\T�Q FL%7����'HbH�c	�<�R�����-xz���'��EE�p�����̆2�(y��'-�{VmJ�l�̘d�+$�@�i�'��P#�قI��T �(�8�'��U���ڞ�I�.��J&"�p�'����O�c�X4��r��b�'��P�φ%"�ْ6ˁ����'_��ÈOl�29(�{fDa�'�J�ub@�
�Ͳ�G�o\�k	�'��Y�� �E�����~�T��	�'���S�$�=�"Q; )�o[�		�'� �b�g��xr�F �*xI�'G���6a�!t��qF�4�)�'���"Ȭ~:"�ieCj�b�'S2���K�J*>�Pa�5H8�	��� J���,A%K�Cd���4g�|"O��"��ȇ|ל-S�f�-Lx��"OH`k&&I+o:�H@�X�?����"O���%��^�`�ā)fZ�@�"O���E헱UQP!hC�(P��B�"O@���E��@sDT�?Dn��"O�J4.G��uт�`���"O��Ha�̈X� \�w �xr�"Onm��2�AA��!���q"O����T�!c ���ś_50"O��W���'��<�h��h�qy�"O�5e-ՍsbL�2�P�|Ɗ�r�"O�0aabЯb_|��b�����-@�"O<�ad��5՘Q�g�Q�L��"O�a���7鸘Y5�b��r�"Otsr��+*��2�iҰk��	�A"O�l�3,>;ZN$0!KR+|>0��$"O�	2��)%|��3I�?DlE0"OĔ� ��0_hhE)�z�n9�"OvT�fQMt�@�0�*��#"O�qI��U;ą3!I�dځ�"O���E���*�`��_Tq�8!�"O.�����5zI��힪:f�A"OlѫP."k������tW�h)�"O�HX��a�����A��Pae"O�d�aĄVF����b�N�"O��w��^�тN�H�(���"O8�%+��Xlu�v�ǲ6�x�"O�X1ҏU������ٗI3Z��F"O!�%���Fl 1Ϯy�
p&"O�qfF�2��P�p�۞;�ڬ+�"O�XӶ�f���� �f����"O�q�`�=�Г�!	�ivƨ�7"O���֌Κou���`g�COE��"O�D����%X��R���7��,jt"O����/R�f4�⢃"`\�M!�"O~@���P�"Й����*QN�ȷ"O񪐩ɔL�~0 1:'�Դ*3"OL�R'�)Ъ� ��җ{�>0��"O���ߚ<V>�R��;N��"O�%�@e��U����X1P�p�4"O�	����k8��F%^"'�137"O��3��-e��J���4S�"O=�A	�1f&\-#��u��!�#"OX���!	.A��9ՂAR�:I��"O�-H��U�1K"|�8HR"O�ERpc"=9ص2�XM�HQA�"OpD�sN�	y��S�F�HӔ)
�"O P����%�N}���#�Nȱ"OZ�P@��fl�	zE��"Ox��t�a��\2�
P=a'xE�"O@[&a� �jx�Ʃ]�J9h˱"O@�;��ԩq� �"i�6 �"O�`����� R�ݬm�=��"OTD@0&��q<����B46�ڑ"O�x2���m�e� �#F��Z4"O���3G�#n�.�p���
��"�"O�4Y�c��i�D��-�K���Yf"O|��W]���xWg`�2�C0�ybOɖ5ބ\��-+a' ���	�y2'��vp�TG@�kkι�t���y��<s��d�� ԩg*H�)�#/�yR�P�rn�z$j��[�R�b���y�I{ㄥ9�ꁉS��0{���y
� �<aG�[L-|ljUo�v�Hb7"O���i�
/[�T�ÿ`F�p`"OJdh�F =K�%$�֭tQ.0�C"O���B�q�uA�#۱/��*%"O�aZ%��4i�D�����5���"O�AA&�B �1���8�  ��"Otq�5��R�U��N]�%Q�<I@,�:
$��`�	������RV�<9ԣ� @  ��   w
  g  �  �  �&  �/  �:  (F  �Q  ]  h  ^r  �{  '�  F�  ��  M�  }�  ��  ��  ��  �  J�  ��  ��  k�  ��  ��  ;�  ��  ��  @ � � / � �% , Z2 �8 �? �E \L LS �Y �a �k �r �z ^� �� Ē � x� Z�  tX�R흱I�8��t#E*��ŋ�4�f���(R� e�'h�Y1�/O�|ڲb�؟�*vB��L�VQ�E�ړ�JQC�D��X+�𤊀�sh���	Ԝ����vfٖ�uw-ځ_��t�H57Y�T�PH#�E��H+3�⨓�o�W�0aQD`[%3��� VI��/�,`�СW�u|ם�(�ؤ����d8s�>;�؄:d�ݾD4���b���Bφ��?i���0t����7%�K�"�BB�'���'�R}D���n=�ȥ�b�?6�'��,���|����?��b� �����?��=7n\B�%^�_��(p6_�?)��䓉?���S��'	�d�0>�8��̙��:Uy�nݳ5!�D�B]��xJe�ԓTo��V�"ʗ0Y_J�a������OMBi��,�X�x+�O�Eyg��9R֘*�LJ(:6�X�Q�'"�'�b�'�2�'HR�����j�pQaWk��JRT�������u�j�o���M{ V�8BݴG��%w���mZ���p�!��3�����;�TY�As�'�^�b#�3�0�WNt"Hs��a��X�����tW~i�1���M#3�i�P7-�t�;�d�F�/Bt��D�*����P2����i�̨�`
ć6ضJB�H�{\��h���ZL`Fk�m�!�M˔� >C$PE��A�F�@ ђ���v�.�s i�<P*v�i�~7�D�����u(UIE�$@@�U�5!��
��-��N�>�	�i����[b��s�$��+P��M±i��6��(~��Ah_9@����'S�Y�f��m�����h�/�� !�O*lȁi�(���2.�72��m�Of���#<]��j��N�T	�R�Ĳ,�:�ӥ���Ms�i��6-���IV0V2Lp���+m�f���S.���D�W�n9ZT0��єC��&�0|�fB 6"F�j1��x�4B�	3f6��4�D�rR|�7&̩\P�B�ɣ%���v�̃i�(�7��;��B�I�5�ZhXa�ڷ9����B�	/J��y�CO�m^��SM�,a���=q5d�^�OD���a�=�`��@�{A�tZ�'����b�b	��)ul�n����'K�L�3�;a�Y+$�"7ʍp	�'Z�Y���+��Q�fQ5�ܠ��'��M�!hB�N�[D��2�j���'�m$ �.P�l�A%�?�P`���>�Ex��I2C�&������2��5���]�~C���<�s�fߚM���BF31TC�8[/>�R�k֟��tP��W�W�B䉐�i8�N^(��F��[?�C�ɛlX,��a6�t��@K�==�C��T6�\�ĬN�"��06���EBtE��ɒ|'�dpf(�(Z�L(5ɈAw�B�I%qx6p�JV��-&��q��C�	�KuR;�6.)�3�j�
FxC�	�(��8��av�ro�_jC�	�['2�p�H�l!�M`��͕	VF����a_��-?iq�&��s" �*�|�؅�l�����Kv�Ȧ�>��Ն:LzYh�m�:�^�(�+}�� !�L&��l���>�ǣ��O~��"�t=6��fT�x��/�Or���O���ǌ_<���@KJNZ�a��A���ʓ�?����i��M�p(3�[Aa�Pp�Fɽ58�r��Or�)���e�Ƅ��nF����R��',�	 V���4�?������#J�D�J�R���%'�f}��j����$�O�P�!	��$c��g��ؼj����j*}��R'%�I�,7,\ q��S(��T���<�8ܒ�c6��	z.=�I۟�'?e�|��f�Y��0� o%�-��`�Il���3t��"J�>�����㍒N�?AU���>D�a�D�GP:���>�ҀnƟ���ҟ<:��їn�9�	ܟ���矼�;+�Z���#�$tB���5��O�nQ��{Ġ�$d��YÅŞS��'��hG%\�r@H$W��p⁕�S���F/@}p(��	.r�$X�&ԭ&9�n�8cw� b��%�����3�� 1��O�c>��O��� �����XQ���+v��4�8D�XP7�?IQ�����t�y!��<���i>���@yr��N��`�� �3(H`����v�|���'a|�o&}^�%�p�	�4$��Q��~@L�2�'6������df�A�P�S	���2'�o!�'͠(hF�_�` �g��z�|a��C?�?��'ߊ�ka��'."��@�^aV�K�'&Bd�R��
vT�5�Č�<ԓK>aºi�'OH��'�		(�pRQ��.��':w3���D�H��� ()��LI�wbi��I��#��B�'	�h�����:�#�cX"
����wL�+�ax����?I���?9�pX"T�%��V{ Ȓ$�fr��.O|��0�)�';�����L������dҮs�l\��	��?1V͊�o�n�S��+h��j��Οԗ'�(@�+u�~���OL�'D�~|K�s�4(�'"CЭ��k�*gl$����?��כ�#�� SN�!��H)t=X�'��ɉ�8i���#to>� ���.t��3p��oZ�!�@�y!���}��'] x/��x�Og���tΖ7���A*F�M�\�)�O\Y!�'�Ғ�$��ĮtzD8��k�
Nl��	O��'��'�(�(�F��d��:eE͞�:�{��D�d�O���B�p��tE�%�y�b\�H�	��$ oØ]�p��I��IƟLͻ ��3�ƒ�"ՎB$��v|,�)��c�AQmV�Q���C���E�'fӉ'ՈȢ��Z�l���B
C�Qݶ<�3���]vѫ� Z��.xPu-�	8�@����@W�'�N����Ҭ�(=�}��b�8""�'��#����Y�8��#�x��Gg�&i���jF9e��ȓX�4���̝:����b����'�#=�'�?I-O��'+�q��0�+��33�S��P�٠��O����O��ۺ[���?�O��8*2vc��@iY Өb��N6�x �D�� ��$.�����xn���'�ƈx�!ET�z�W�Ѫ>ѣC���?��䓴?!���'��	���f䩅�.2��r6"O��s"<$��D�W`�|,t�4�|��y�Z���<qW��<Iɟr�ꔄ���LEk�+3**D���'����o�*�(�扝[�`q�fj_���[� ����6h�qO�Dۇ�Úi���j�&Z7�%Se�'�L���?�Ol���	�#����J����'/"�'��OQ>��l��!�܀I�#>N��B�4�O�\�	�@�$XZ��$$b P����"�	�a~V"|:�w��!B�G���]�ȇdϘa�
�'�0ӈ��̮ő�dU�a�$���'�` �wL׸;U( ��;_����'Vv�����.�0a��W�]e�@�'-,X�"��Y�=q����O�8q�'r!Yf'��z����Bgd���Z�8�Ex��i	�=5䬸�O�e�d	�&�\C�IP���)$=�`eHE�S�jnB�$3<򕒲�A� My�̦9�.B�	�/��P�+�T�yrg��B��5s�J�'�D��"	^K
�C�ɌK����S&<l��UzgX���NЅ��E��� cj��4�z����C䉞5�du�#G)nI�&@Z�.�B�I65��e���ͥM��
6�:zB�I2x��[WJ�<u�:�撒y��C�%$�*� ���H=ɻ$aO�L{\����93����3|R�*��¹l����y�!�$^
:Ҧ,��ʝ/;f`��F�;7�!��G�T���/.D
f
v�!�ؗ[�� �c��V��%��O>!�d��3zQ ��v�x���3N!�	�5����4�@3G�KALў̒��2�w�l��"	��1�T��F�]�~��ȓ�n�3�e9�~����3_���ȓ*X��c�
\#9J��W-�;"v��}q�1
Q�.DH��BgH�X���f��bK|����س&] P��e�y��#;�ࠂ�n����I���"<E��̥ cL�G��!&<�[Y�!��Y�t�@��p���� Kj�!�$��IsdǑ0z]t4p%�&1�!��P�F8�cNDNJ�]"��B�!��Ao9nu{���7^� (��S�?!�Dşh ��8=Pb�15E8��ɘ%
���AVX��1�ҕP���$^9{!�� �=�G�ál�R���j�\1�h�G"Op���B�+F6�*�i��&p��!"O�1�i�9W����[���%p�"O�%	����h����Ǟ�2J!0w�'�����'VХB�ȱ}�l�S��W�!��	�'�<�g�*�<$�산�ƹ��' ���eۄ�(���V4��
�'(�hӬD�4�b	8�(�����
�'g����h���y@G�Ll�(	�'~��t&1=��[���G1D����I;`�Q?��a�O�����lN�h_���0�3D��"�A ��:�kBI�
��x���2D���MH\�,H0E�T.;�jd��0D�D����"Ky�L��`��9#D� �G$�t.��è� �ap�I$D��Z�40����Q�Z*옸'��O>����)�'0�*�Q!�w2r�Qd��baKLT�<y�@��a�uA�oP�,���Ҵ�K�<�Ū�5���Yu���6mr���H�<A[	p��X���@Q:�;V"�!�0o�\�����Y���A(�!�$��Eح���؉ Gd<�c(D��ɼ�|����4RH��v/U8$��4`�I��D\!򤈋�^}����ea���0(D�R<!�D���(3a�ʱ|�����Ȁ� !�d�3G�̙,D�F� �J�r�!�d�s���DC�e~& q6��}����~���,�2u*� 26�8����y���E3|�2�-@�&y�!Q1+���y� ��(z9�����!b����[��yb-T�}���A�j}:�p�ϧ�y�hZ�~19F�
id����mů�y�nŒD��f�)`� l�&��hO�Q�F��_\Ppq��7)�VY�u�I� 8�C�I�t^�9";#�C��7�C�	0o��7LW	�`D�B5\OHB䉵5;�Q#Bg[�*��B���C�NC�I�/�����a�6O����dB$ �lC�I cA♪��H+�pH��o�;Z���Ae'�"~�W,��2�U��O6�2Ȣ��Z�y���?����p�
�Ά5Q�D%�yrA	J(�Q�c����U@�y�K�!��h�U@�w�$�+b�[��y��Rd�g&�!m�fTJ1�H��yBEP����3U�Hd}���p���$�>\��|b�('�`ӣ�1���r�����y�
��r�&؃��W�$����G'�#�yB
�=`\YS��;i[���6O؛�y��o	Y�B�h��5*��R�y��S 0�MҔA��Z����n���>���e?-����]�F�^I�/;Ni�ȓo[ ��6�/P���T�Ȭg�4��P�BA�h��'�^��'�]�lb��ȓ	��=���Sy���BY-��م�D~��U��Fl���ޭ
L�ȓ%\�yQ�L#x%�W�N,d��<G{��(���R�eN)LNt�{�cR�ld�g"O�|�n�/|~h���Ȭ#��H�@"O����WqPd��� ^8�+R"O��Rt���o"d���U�4ư$��"O
���H�[L8��O�!y�"OB!�7� aeDŋ_HԐ	R�'�M����S�~�e��9���0���긅��<� Q`��;} <X4��5qL���S�? �I҃�z���Q ƍ:���"O�h��k
\����%-Ӛ�:"O SBM� ~Dj�+ۥ�Fqɐ"O��R*͑�jm�1j��$��8�^��QB�9�O�)qU���j���Q L9�!�J�V^����u��s�|A!��Y r��r� -9X�b҉�8A]!�$R�/�j#�Iה[�*��ڈ/�!�$� P���M�6,.�h!d��}��ļ�~�˪6�l���@����y2��A�d�5�[�s$�����y�/�~V"�Hա�4;�HkƄ�y���1I�Li���!0x4e�4� �y�#ǈ�P�21 !�*�JW!��yR�ZR�8���J�u�KV���hOp�Z!�ӑy�v��2��\��aZe�V�Y��C䉹6gB��7�S��D/ߕk��C䉈Y��kG�Θk^�1*�&ߨA�ZB�8�6�p��V�jގ�A�]:UIbC�I>�8�ɢES� ȜU�ѡ]O�ZC䉪�$'&��!ӄ����=b�Ğ��"~J �
�������p��]�/��y�)�4ۤy�Ck (c"��R�-M5�y��.�xUhGʟ1)��@0',��y�e�xN�Q�e T�;F���ϒ=�y�ȋ+%�Y7� 6v�Ĉv��5�yBBY?rH����'W�ļpf�����Qa�|b$�^b��ϖ�#�䐲�	Ɵ�y�Dd���I�!� 	{�	��y�����KE��)�i���[��y�/17t�H����
�ʉ%�yrA�z㐕�B��_��3@i����>ɷ�GY?a�d!W��uBSF�;� �RU�<�T	%ԕ��iWk6u9���{�<�Rn�*n�j|a�&]�';ZY�1�z�<�W@���B�H%g�v�|�<���V�0̸aAO
@V��pU˄o�<�ڜmU�!��J�1�m��Zk�'Rx�Q���I�h���<]�h�W��<�!�Q�R�V�H�+�7s"
���Ö\�!����޴�t*��
B �4�K24�!��,v]��g�?	��Y2 �#9�!��7	JN�ŭ�P'�}��,�u�!��
� m.�C�\´Y�l@�,y"	���O?�QӎM�r��YF(��l�0�BTc�X�<9B� ��+���I`2U:��_@�<	�-YL��Zd%�	�hM
d#w�<ID��%rz�a览
\J���a��u�<i�(<�y`�c�V�bْ��t�<qdF�E����,\�}&:���lDfy�A�p>aq�I�3���Y@U;2�nܘ`�m�<���	4�ճ�b��8vL!"�t�<�U�!im*�"�/F�K�"%QP��m�<����qi�\#d�G�j�p��u��r�<�C]�
	"��&G�O�N�`��kx�p�n��س�C�E�n=9T�H�i�Ry�3�2D��b�`
L���aaB��0�9��2D�P��C1x �YTKB�s�q3�/D�D��b��(��Ѳ��C����w�"D�$Ȧ��Aj cg\'���A�,D��`�F�SwL(�F�$����D&ړf�f@F�ԥ� Kʼ�p��̟2I�(�T���yr�ش}��%�Ӿ"���K�,�%�y�&��m�"D��O�
�ڳO&�y
� *��'"�O�^Iҥ Wo(8�"OP��R�+���#�#�!zZ�,��"O���u�-6�Gc9+8�A�'�,�����(=b��T�� ?є�sQH������mL���$
�mo����=	m@��ȓNnNh�#�
f<.P%���]P����?�`�h�Y6$���(�5򄽅�Z߾���i�#Z(Ma�^1=�|y�ȓ*�$�a��EK:P{B�,j=�q�'���N�h@��&�\��h�h�x{t��m*�Z@&
%��(hU��s�*��ȓ���g֊~C�=�7d�ErR��ȓ�Ĕ�F�Όbn�0b�nD�5�@d��S>�hsǦ�8s|���R2]�J����"P��I�?���"�b�hS���Q�B�ɛ0�X䈥��\��`�Į�nS�C��>����������
U�[��C�ɨ
����P8洨x$�2fC��(R���`����Y!���zo@C�	;}6L@����ܸ��(��	�D�=�6�@r�O-���GJ�(s�M��Ʉ�X�|z�'^�!#�k�+Y|V��OעH��,�
�'`2�`�#Ȣ���&��*�B	��'jr��d$S��6-�K$8��'���&I�4298�.��q>�M�'!(tZAi��(�(Y�ƀ<Z��z�jk��Ex��iEj@m�&*�
�� �D�G3�nC�ɜ����vN�|Ԅ��n��u
bC��9v))j��D8/�<|��`�F��B�I1
b�hb�5%$䢄K�k+lB��2{�@�`���G�(	�o�1	.B㉉K`
����93�ti�M?���cc�_�-�Jh0#G\�"����?1�6bMw�6\$�?�w��y#�)L�VFax������c0U����?���y�V����^-i XU�q��>ͧ�"U�"(��Lk&� u�¥K`�G|�E_9^8إ�o�7%ά�0p����6N
�M�W��%(`��V�ɇ/Wx��O�c>�02f/�"��fB[;�F�a�f�<����0�uc@�:hz(��!(Tم�I���$;�]�֌ğ�j�:��>F,削S�T�I	8����g?���^V6P!%��LaV4��$�<��N�e>�D�d**!�����iO?x7���(�7�֭�ả�
�'��9gAٓa���BҵD�?=�/"ɶ�kFƕ!�ek�,Y7�y�۸�?�������䜟P��Y	`�e)��X�Ov<��@�&D�X��`؋p=X,a�d�

ԩ�F ړ~)�?	#/�=�
�:�EپN��+Q#@�<��?��g�'�"��X��+�+�F10�ӑ�Z��yRcTQ��A�IM	B1�� ��(�y�c�hj2쓱 A�.�ǋ
�y�o_�}�0��tBG�?�l�As)ѿ�yk˶3	��A��F"	6��Kr�J)�yB��p"V�h��J�UEi�q��"�?�Ѝ�v��0����=�%�q�	H��ԩ>D�h[Fk�0y�+��͓PzZA�sf;D����BC�%�4�p�Y�f�`���5D��1�Ŝi]ʘA��2�*a��>D��KA���l��DA82. ��G�>|O�y��>�jϟ2Wư��P�xv�[w*�x�<�$΄(iC8�I���,T� �d��l�<���C	��	0��0&�i�<�"�	Kl�e�PiB
P�nH8�e�<	 �3#��u�N&�7Od�<2N �1����(̋d�����v�*��mFxJ?#��7Ұ`�׷V�|ey�;D���rEc�HFKU�xw:�Jp9D��pN��b�0�@� "XF�y��8D�� �1��e����+���P��5"Ojq��U,<�����!iH{S"O!�3cAzn�\����v�Ա�T�Ν�Ot�}�T�0�!�F�\PIR נp���`E��B�h�]���Go�p���c���M��s�����؄y�¡�ȓAm�5�v��esT��僟?�~l�ȓu�����\	AfX�`h�I����ȓF���Y���J�icq���b���"J�����v�|qʕ`ވ%��	�F��� �!�^�KBxh��F��&5�qN��?�!� 9e�N����
<W��I����!�D�:���RCH�w�|A�%��i�!�D̸d�:Ly'G���>`����џ02R�y���|B�HݛR��M�p �O�4`�a�b�'*�%"�ld�O�PE�"��M��ii���Z ��$Z7y��p��i��
�NQK��#D8q��źU�HP�O��D'�	#f�~x�%`��$�
�8v��&�����O��"~�1 ͒'�@�C7�YC4h���GI���>y7X�Իgƞ$5��0�A���G�҄Y�h�<���?����Oh���!�&��K<F�0T��W#�f��� �Y� xS�̈́ �*���EK� ��	�?�ݴ�ēBLc>�A���"Kg�M�Q��ѷ#9?!��O��G�>��y��L��MSצ��)Ϥ<�ъ4'�m�4&2?iԚ>��e�d�d�vⓐچpF��.g��
�#U+K�Q�>i�O�}�&cVq�G]7l��A&B<w�:��bF�X�$B��t��t���(�:F�;*�\���+�h�z�B.c��ܚ�D�D�N�����%��ʱF�7�$�����I�p�h�'�V7mJ�
�y
����x�C�|�ɬ#��'Y�#R2Ă�a�Lm;u��8?rfyxg�� ����3��S��'��ȑ�OF�#�ʊK��b�	\4Bx��e���ʤ�q���'VL�P�'�1�^t�#J����B��Y�t��'��<�^����9O>�H��Ol�e�\sȜ)hV��:��ѡ�'�҉��	Hm,��#FP�!(V��l+�B�1	Z����9�|a��C�
�R7��OH�O������|n��4a�Ѫ�q�i� ��L�����hO�S�Vbބ�r��!6`�%k�$(6C�$9��'߿\ʄqPN <��B�9�����-n��$�߁�.B�I�f��-E �8�!�2h��Hi�"Oܠ�.�u����E"|T��"O��G�N8�|�Qe[�U��X$"O��2���4&U��� $f����"O(���K�H�h�j�Θ`V`�V"O���Α.����`L_!<p�"O���n��'�Rd�tk@�X����"O��i�ݘwQФ��JJ�T,����	ß��������Ο�����!�\l��ņ)VW`��f��M���?I��?���?I��?����?�#dC	�ZMhу�=x�{�aI.͛��'P2�'H��'&��'5��'-ң��u(Y�2S�v�Ґ��c�26��Ol���O���O��d�On���O��d�%��X"u���2]���R!��8+�lǟ4�����	ܟ�����<�	��	Ka�k���c��JE���ߴ�?����?����?q���?I���?	�imPh��/]�O����g҇|�8q�iz��'M��'Rr�'�2�'�'4��R��ޯ[�.��@jK�>`l���l�H���O��$�O����O��d�O��d�O�٣��<BPI:F���W;ԅ�T
���)�I�<���L��ݟ����������y�#�+�)��ֻ&�|�	��M����?A��?i���?����?	��?1�`Q�r2�$�P�J
tU���7 ])l����'��'�2�'���'���'�BM9|?"���<cFj �*I�G��6��O��$�OT���OR�d�O��$�O���EMV  Qi�]&6s�
�V4L�m����	���Iן��I֟���ӟ`�� _�-���N=!���ER�j��Q��4��D�O�˓�����A�hڤ:����)\�f�Z=*p�t�<��F�D<���M�'[���Viȍ_l����c᠌��?���y�U�'?�WI��a��X�|	��-Z�o�������>V`���<�v�'	^F{�O��d],!�k����5|��E�n�R��$�P�ܴ�)�<		� ��H����˵��������t}��'��0O��'r��ᵂ�_��Q�ߗ`�쁕'/R��\a�5��O� �?a)l�P����
�Px�$푷o^�C�<I)O��$*�g?Av��G��tYG��"&�	#(��4�޴f��Y�'��7�)�i>1��M֓�Nى��RW�$M�4k��<��͟@�ɛV9��ou~�1�(��S��S��
c��S�Е{��9�DEK�',RW�X�|�P$W�E$�z��T�x[�l��V]yrkz��m�P�D0��;R��p	�f�ҘQ�!�5�Jl�O����O
�W�O���(ebl�$�0v�S�$ϔe�f[B%�d��O��č6�?��+5��<A5� 4��6l�[��5�l��?i��?���?y�����eXh��8�nԹ�����ʷB.���(	蟤;�4��'�ꓯ?��y2�Ɩ]��8R�T�Skf`�ZBDl��4��$��G=R����l$��x��
.D�*���
Yj� ���:}�@�d�OD�$�O����O��:§<�9���B$	��1��/�pTE���p�	��M�LĪ��DΦ��<���@�}YԌKԢ�:��c���^��ڟ��	ޟ�xB�Цm�uW�@|��TE�/��㠋,��Ї�'_�&����M���?���(pHy��4F��6,�:X�и��?�(O1oړH�>Y�'���?}0�FV"@��]8PN�2X4����Or���O}��'���|J?�ɐ�L�p�`.�9s�r=AF��(Q���R��	�r˓�����O2 �O>���=y�c�h�m^�p�qŅ���?Iǳi2���"�A#*�Q+�� -&t�����*��	0�M�2̠>���NH�Z���*����n�vd�����?�C�?�M��OP}��)���T�?�2���y��q@�)�1����O�˓�?1���?y��?������ƽ.B�ap���;�ޅ`�,S17��6�f˓�?QM~R���&:O��I���e�@՘GG����¦�'�Ҟ|����L=;����O�lJ�h_�yVl݊tEK�y��i"�'����g��,�ǟ|"T����Ο���H[�}ki�3�)��� &��՟��Iܟ0��Cyr�t��œ���O�D�O�(�$���,�ĦD�f��}i�(�����$�O���%�$ox��W��u�6Y�v�9�����R�IP-g��	��d����$8O��i�!�~���O�$���6�'?r�'�b�'Z�>�͓�H�����5H�V�k�MK����	��M��
�?����V�|�O��T�kHp{2���{��
?s���'���'�����i��	:%�^5��ߟ ���H�2z^�+4	\?j�aaI:�d�<���?y���?����?TcJ�r����O;�
��ADO���\צ�R Oy��'��O�ች#��oT+P6���L��H��ꓸ?����S�'6H\�d��8,��B%뇙{"t�,L=�M3�S������de�.�$�<���2����
M��3w���?���?���?�����d�����J�<�q���w�0js�ô%EƉҶlM��Haش���?1UR����� Γ]m��r,
�?#�0�p�W� ��4������'���FWZ�H~ʛwN��D���0� ܯ	t��Y��?���?����?�����?�S��JX��C�GM�$Ga�?Z&L���?YŻi�(����'���'�2[�XBlФQ �`�	i!��0�\t��韔�	�(��L��5̓�?���� N���QdB�;�r4�3�̪pp�$�j�O4t�K>�-O�	�O��d�OJ�K�KN2k��5���eL���,;��'^�I��M#a��?����?9Ο�D�VO��V�0�x� �"8�6!�_����O��d�O�O�3�rA���J!PTư>X�(:�,דpČ �APy��O_�a��u	�'[�0G���0 �`�nA�/��N^B�'�b�'���'���Ӈ�'R���M�d�	352�J�
�*����`雏;��(��?��?�+O�$�<���rk�e��#9�FEb��D�=���?�eOˊ�M3�'��G7r%��S�����"�p�+oL�mfb]�R�k�i���ß��������͟��o�DK����	��cѳOA��� F��6/^�!���8$?Q���M{�'�Zd�� �(6{��Jdf��lz x"��?qK>!K~za�/�M��'sd̰��N���cs��4D�D�P��+�h�����'�̔'���'O�A�jր".��2NP�iϜ	+��'���'�r]�${�4m��i�-OD�_�F8�G�ɧvWn9{D��Bx����O����O~�O8���"G/�y�RM�O
�����<Y�O5y��T�ݴ��4����'���7J$Y�7U��d�Q'�B�'�B�'����<	�[<$D�T�<&���F��� �ش����?I��i��O��X*hBA��Y+m�i9%B��$�O����O��	��g��nZ&�h�A��]�@mn�Zt��k	�帰�$辒O���?���?9��?���J�.|;��@4U�\ȉv�_�T�J**O<IoZ�����П(��h�ПH�M� O�R�2��17�6�v퓊����OH�d8���Ы@�� ��:JK��wb�p�Xq!��
	FZʓp vu��e�O0!K>�-Oʠ��ĳ:�V0񧐮U�`5:�
�O����O����O����<Ig�in�Q�5O� "-�򂐉r�� M��f���'�Z7#�d�OF�'R2�'9���h��
b� 0$�h|�bIҨs�,902�i'��%I�Ρ�Aٟ|��~�]=p��="C���-8�a]0`p���O|���Op��OH��%§o��8f��fI������-g. �'<"iy��c��OP����M&��Hf�вB��U�ˆS)r@0�e�~��֟@�	���������'��9�y@����ݗ&����MV�x��`��������Or���O>��23tha�&��3����S�H��$�Od�~
�vk�=j�'�Ҝ?E�gYDx
%jE�.І��G�<	A[��	�l$��O|�q�&đ,�z��@��V�R�9Ǉ�Gjr�p'�FE~b�O����I�
�'�RA��)ؠJ��rÍ�!��1V�'��7��V6b�q5�UY��t���k)�]Bu��<�Ƹip�O���'�B'ںR�l!���9y�B��L"a��'�d�e�i���&[ȸ�r!ޟP�'f��,h�,p�~)�wOЉ=�Ό��By��'��'R2�'���?�P��ty�4���
e�� ����9���^y"�'��O\�/c��~�P�`!�R8@��!�M%d���Ov�O��,�R7b~��	�30���&e� ���%�>k{�����]Жej�X��O�˓�?��c��0c�2$�=�2�\�}�U����?q��?�-O��m�=RM�����	�W�j�Q�M�]��X8�Ϊ5 �?AT���I�P$��ц8�<�҄`�&(<���}y�K�	>�`�i�x��8x:�'���X�PQZ������L%q��$�OZ���Oh��<ڧ�yB�ļt�$��aP�I|����K�?�V�i��E�t�'XҥiӺ�O�)���}*F
��M�G� ����c�O��D�O4�$5*YZ6M8?�������g��
�̈=]��K��,��p���/��<����?y��?����?�rLEX��ہ+B�k:(a�W������](��Iy��':�O�BD�$�	�#�׳{���Uf�(=���?�����S�';����*��\���T�v!�CG�Ms�U��2���<��"���<�@	��i�iZ�NѵS2| �Ǎ���=��i1F�18OvЫ���|�>�y�&��`P`�3��'U�7�9�����$�O��Da�t����;~��h�si��uU4��a'�r�86�>?����t\8��D����DKV�S`�q�׈�$,��C��P�	���ܟ �	���F��k��U pHr�ΦI7��v�U�?i��?��i$�����'���o�Nc�H�dM�"(�\�{�/�-%� ���=�$�O ���Or�2��~�2�ӺKf�\�m�xܲ��H.I�������^��]��nX�O���?q��?)�4�b�*P����안�̴5���q���?)*O� o�R�v9�'=��?���� ZG���UB�	l�a'��O��DE}b�'�B�|J?Y�-� QK~٘Վ$Vn�a�%�]ќ�'�a�q�'o��E^y?�H>�" ��%e����d����	g����?���?	��?Q����ɢ<��i�z�1�L����(A���>�i��j��S���'�>7M#���O�Q�'o���-A'v�X���@�δ�R�2@���',���g�i8���OL�򰀆��B祿<9�"P��j4`0��7t8�u&�2�?�(O��$�O��D�O���O��'=��e�g':M�*}A���%l�D)2ٴL�� j/O6��7���O��o��<!�`�gU`��c,�,e���D�\ɟ��Z�Ii�2�" 4��z�|��oUf�̊���A-l�䗊 �|�@�'U�'��	՟���:C����֔/ơAU-ʌU��$�	��	ɟ��'��7틱>�@��?!%���L���	( �ath���䓂?��Z����ԟ$�ĸ�#V�C�
�G�c���K�
cy2@��МÕ%Y(��O�Ԁ��*���H(2���D�SV��<Kg�ñ7<"�'i��'r�S�<�#i3(t���d��m�w����ٴB{dx��?�a�ikɧ�$�Ok��xF�O||�L)r�	#�h���'4��'R�����֝5�t���g|8� ����e��ƕg��d0�|�^���̟����8��ß� ��#�,�E���7¸��ˉIy�g}�L@8��<��䧖?��I�3�B���P�p��C4��	����ID�)�S�h4�y��	Y�-���bA`D?@�X�G����**O��d����~��'��	Dy� «c,|�pa�'}��aG&�4���'P�'#��',�	��M�)��?Q�X2*����$�+v��TrW����?�½i��O���'L��'��B+I�<�Q�J^���8ջ)�0�W�i��I4Tۦ@���Ozq����%|F(�"3�ǭ#��RQݥVp���O���Od��O���#§(�|��v�ۨa��8�EY�l�Α�'��a{Ӫ��d.�Ot����u$��hp(�l�RT�^B�P:q�H�Iǟ�	ȟ̻1	�Y�'!K���9����ʑ]bꄪ�G���������O����O��d�(}) ��3dїgG��+0HF=C�p���Oh���N*@�I����O�X��AǴs����qgE�}�h���?�`Z���IݟH&��O����p��m� �
�f���J������n�CJ���� (��@�@�O����	�.kڐx���G}B͠g��O���Ox���O��$ʓ[�f� �u��IRY|��1pO	�P(x%���\��	>�M��O�>Y�l�h�r�H�P?,���K��\t2��?�b_��M��O��3������?5@P�D1���pc�5���pD��O��?!��?���?����i]�4^6<E�٧mf�$��ML�4�n7��=_����O��D<�9O�!m��<q� �?y�d�`&��ʄ�����l�It��~�7��n�T?Aq�<7��a����4�����sӫ�"���9�$�<�'�?a' !(�x;c���c�$�z��H1�?Q��?�����֦�ʒh fyB�'��� �%UE4`��hI�c�9���|�'7B��?)��� @8����*��D��܀Cz*�*O�D*M�Y26-LD��:��k� ����3fzp�eb�-B)������O�D�O����O��}��'�U+�I�T�T0�"U`��X�-ƛL
c"�'df6-*���?E�,���D ���ċpV�5�`�ӟ��	����	�DL,)o�S~�"��w�&��'w��ř3���M9p(«�$u��{I>1*O\���Or�D�O��D�O��0�-�	 Y,��1J�$G���	���<��iR$,���'���'��O�"n�v.)��ٛw�!��<;vb��?����Ş&RdU!`�ݢg=̘!�r�dE�&��<�MkwX��'/
�x��9�d�<yv��5>D� ��Ni���QDaÆ�?A���?	���?������馵Y�A�ퟸ(aʙ�d{���A�I�rq�`Yޟ�ߴ��'r���?����yr I�_�t�;�nJ�/�b���E�1):r�4��duC�`�O��Op�n�H0Lhr���gR� j5���}>�'"2�'���'
�����'�6���մ$��-�Wd��1w>�kE�܇P���'t�6mY6C�`���O�oZ\�	%r��պj4CUX��r���-�r�$���	ן�y�d�HwӔ�ٟ��z��I	�珸,U ���^e��#Q!�՟��|bQ�tDx�TV�	9�K΍ ���+��'�&7�N�R,R˓�?1Ο�X��^@5�0C�����h�T�� �O���O��O�'w��8��CM�dJ&x�!�	g٤q�NϨf��mZ��D�h1�'�'���Y��d�L�D��R�sg�'�&7���,��t��%�1I�(U2��C	 N6�ᢨ�<���i�O0U�'�R�Xr���c�<�$�3ec�v-R�'���AT�i��	�c#숰Gߟ��AU�x2�+ɱF�T�a��$�tM��gy��'hr�'�2�'eB�?� G�	�X<%¶AGcV,;�ڦ�5n�����ɟ�'?�	��M�'w�]��^�zX�X;��?eQ\-���?�O>�K~r�� 7�Mk�'v��S��t�R	a0�7Bֵ��d T����O�qcӓ�lؠ�C�)�n�{�E^�i�ڄ�ȓk���#G�R4 �<<��CҬK�����R���	��pm����1F����5�o��	��խl�$��5nY�%�������*n���
G.*@U����$b� �aAoӈ4Q�Z��TRgǟ.dPvJ8Y�580̓'���L ���b
j�9�FÚG�X�1`�1.:��&��d	��@C  
J��3D��mf����X#�����'LBH�e盅[��`^*.5�2l`�!B"N#R�6�K�k�?4��q�'��LR��!a�Z<�%k��UP�	H�d��*��D!]�4 ��Kށ���6͎�l�`Dr%�z���h�	M�ptr�9�i0k��@�7O�*� �:��J�5�^�EG�,Q	q��U�d�Co*_��ѴJ�ð���O�!)m��/�UZ��6�H�_���V�]6�`���"R�~ܰ2"yD���i��'W��OvȬ��E�]�(PB�菿��}32�|��'����O �(7
���3��SƔ@*�N��! ��$�<Q�j�:#՛��'m��'���Ⱥ>A�X��Vh�/�
�P4���?����?1f�	��'\1���6��4g�Œ� ��{���'�D�B3{�|���OV�d���l�'�剐e!
�R�g��.!�E��i P|����|�5�?�����'��q[ԦO�o�q��>`;	Az�v�d�Op���8&²E�'n�	ǟ��aD}�b"��Uo$x
3��A.J��?!PkP��?����?�.�Dk6��DФh��?i��N?��X-O��$�O8�d1��) cbQِͱ@,�py��]
�
@K>	��?1����$L;:�j���z.ƈ{��b��D��j}bV����}�I�I�BŃb��>.��$Q7ɤ
ш=���|���p�	���'CR|*v���8��$^���݊É*1Z8��'M�Iџ�$���	џ聍D�<	��Z@�س.�6'�" TlNy��'���'9剿#�pe�O=��%����'M0+�50a�3���'[�'���'�b� �'�	,<�T�h�@Q'��k��9� �d�O���<�Ȇ���i�O���;��\Eʔ0�]�K�Q�E�2���O��$A������h$��P��#H��!�-S������<13Eͷ�V�'��'6�4/�>�� ]*]>����r}�h�)�?����?ic�T���'1���H�LU4@�Z���O�P� ����'F�E��e�����O\���F�$��3NVL��oȾH����C*O����	��\�	�&���<���Du�|��Z�v�R��MJ�\>�@f�i���'���H*�O�)�OR�I�g	�$�T�\�-��q���H�D�OȓOX��<1��?Q�7|L����ueƌ�b�A�J����?�a�]5���4�'��'�� �p���e�� �ɇ�'Z"Y��|B�'w�'G�Y� �I�LK��2/Ǯ�Z �$CA:jf��с�_y��'{2�D�O��ɏqy�$�Ɔ��Z���B�7���Đ��	ޟ�	꟔�'�l�����؛Pk�89�6 �"Cn����Y����П�%�����T�'�$ɻ�BD�ƥQ5��e\�84�|r�'n�	˟X*�c�X���';�ptGW��	�Ĺ+JVI��'6�O���<��j�䆨a>פK����
�cY�7�B�'u��ϟ�DO�O���'+�>�20R�a�.+7n]B�NT wh��7�|��'~�8>ER#<�����(Z&/��'֍{aȃ��?�(OJeY'NR��O���Oz˓_����D��c$"� @iB�x���	Ky��'S��Ԓ�Ԃ�E�2���;lƸK�)�=W�2���C���'��'K��^��'4z��S�^y �Ӡ�\ C�i�/O|��)����Ty��M�	1�n�>m���{6 ��Ms���?��� ���x�Ox�=O��H�0) pf�ɞ\u:h���'���|bV>�	�����˟8��A|7؝hc�ł9���C�Z���ɻ	^��K<ͧ�?O>!��͟��PP[P1�4�6	�p�SH>������?�/O�dBt��q:�Q	nX��bƽr{�|�U��<���?Y���'
��,}E6h�wk��QyV	#r`�$��\)��'6�^���ɋ�r�'.}���C��qZ�5�q���o�m��ퟜ�	c��?i,OȌ�ְ#E��a�κWtM�m)5(��?���?�,O�UzUt�S�����&	�VInf���e{D���Ο(��ay��':�Ƛ�O8�Ƀ��9?ֈ�����;�Y��'vX���ɨ5�b$�O��'��t�����cĉg �U1B�#O�'!S�8	e8XR��H�`�$��U�� �>������ė`��n[�4�'v��b�<1G�T���� !L�hW�dh�� ֟��'RR�'s�OR�O1J	��or� [���]'H���'�h�&h�&���O����t%��$��öF�*1�h��׹c�	���I̟�'���<���v�2	Ӷb[�QT�
�mG�f*��Q�i��'�RɆ?����'��'���'�"ɰ��S�<"dQ��j��Y�X�G�'2R�Pz#�]�����Ο$X�M&�R a�K�Vr�Iz3mޟ$�	�W��dr�O�ʓ�?Q,O��(�X�%ǟ,r�x��ϫ)ؖ���O���7O��D�O��d�Ol��<!�Lڪ�`��aO�Ym��N6aG��_��'�]�������	�G��(�,#aw�s��ͣhk�(��o��'���'CR�'�¦8bp6m�l_� gS�5zR��4�)����O$��O��D�O�ʓ�?ї�
�|��"P+@��q�	�Xm�eI�NÌ�?����?!��?�+OlD�#�[�$7�^M�u�Dyhۖ@�&d�d좡�'F�P���֟��?D@��|:r�y��!��îu>x��ǔ�?	���?Q/O���!FCh�$�'�"�O�v���fF�ʥ��j�Pj�5��S����꟬��a0�z�	�|BD����(ȲG�?����/�ڟܖ'�z�2kg�D���O��䟖��'�H���@�$�H�ڣV1��6�'
r�'?���'�';1�\mI��_r �-���P�|�����'[�)�mx�d�$�O��d�D �'�剸i��0E��]a�(���}��IK4��ӟ��'+��$�A�����fG/�\�c6$�V�*�mݟ���˟DZwoQ���d�<���y�c�	m�r�k� 4x���Cd��<�N>q��GB̧�?����?�6"n�z�gF�6Vv�}נ�?����rm�RW�h�'XrT�lͻ>8� q��A(Et��Be�T�^��'�Tl�'>��'q��'�s����� D��9&�*���կ����[�OHʓ�?I/OJ���OX��H@t�0+N�?�Z8YSE�5�q��2O����O"���O\�D�<���?3_�T˟m��H8��D�t�0����?�.O��<���?I��t�(M�mT��ņ��[��`���V{�Hb��?����?a����dJ�4��O��nI�&�&�3W��S[���������'F�	����I��!�Ov��O�>�J1��w� M�0����=ò�'��'R剎I�P�b������O��i U~���"�5s
�ܑb�r����?���?1���<������m>Q@�*��&��Dy��A/I�Ũ���O��G�
 Y �ig��'Wb�O�b�h�V��L	b����M�pXV1����?)�:Vt���?�.Ohb>i�g���h�z��f�f�����*�O��RtLM���I������?I�O�˓{M� �\�� -m�&�k�VGT�	��`�'�.�D:b�e+���8X�=` (1��mZ�X����$qA�^
����<A��yB)Ơ W�I��ԥz�I@���?9���򤁳<	����D�O��HJ��H;���-n���ƚ�+���O��8T�^h}RX����yyB8���c�,
��A�d�~4���'a��y��'R�'���'��	�s_��9���2*��R�B�0HXB�YC`[#���<I���$�O���O<4Ys�PEj���%�_�\Lљ����R0�<��?�����ă3Z����r�Hn4bw)3o�I�R[�$����H&� ������fh�X� ��� E �o ���P1�,�wY��������ey�ɉ����YPFO�����6pS��Jc��O6��-���O4��$:Y��$=?�@J�3\�)V�H�"��	z�@�ޟ$�I՟p�'ǌ��҉,���O>���WP��q��)��9���	�!힒O����O��G3OB�O��S&-l虗��p�(x�Q  5kq���<IE�cכU>Q�I�?��.O��VcV�=L
� c/T>-X��'�'4��'��(���>��pV\dKʭv�2�pe��z�V�d��R���nZ�0��ʟ,����'�N�������f1k�H'^��D��'��DÃ�'��'��H���4Z��)���+`ڸ@�l�Ao�柴�	۟��O��'��0O��O-�TAi��H�%�,�hF�dV�%��<����?9�Ov:�Qg�"lx�E_�yA�<����?�*R�k\�'0��'��'12��Pn��H���f��>��,B�_��ȕj|���'��'>�O�d:��ED0P� g�߆N��ạ��9c^b����E�I����I�U`Z���ҦUsp|�`O90u��s���p�'���'��Y�У7�����Bͤ=.- ��	�v��; gLq�I���'�(�	���� ���HЩC	*�Ơ�S�����my��'���'��I�+j8!M|bN�a�L�c� ��Q���r��$�?�����?�.�V�y����T��zA@Iu��ғ���?9��?Y/O 9��.�{�ߟ��S._��M*v�P�eb�Cf��.��%����ܟ�c���䟘'���'h����D�W@�[2@�V�>���Py¥��m�^7ͬ|j��*�Z�xC�V	4���;���E pt�`��Ob���OX���F�OV�Oq��9h�# �k��H�KӫCM���D�'Y� ���n�B���Ol�$韄�%���p�`5�e(A����xP,�'eB��	�O��ׁ�<5bH�P�Ҽ:����E��OD�D�O(��ɻ#4N�d4���On�ɑYV��r�ĸ���Z�c�!.�g�	~�Sٟ�����(�cT<-� ��d���C�����U���ɘN��h!L<���?QJ>����90X���#.j:��fC���O����O��$�<w��M�$����5��"�i��"�R|�x�'$�|�'%R�L�&^� � 
�=`X��GC8���y��'FV�d��oX\̧=D�L9fH�#�Li	��A[�u�	֟���Ο0$����Ny"�Ю[X�A���R߂�+L@�t���Uh%��ΟP�I񟐔'^�˄�.��ݝ�~��T/����M�W'�"L�J���OҒOH��+�����%��_�6�bu���]�$��	����	iy��ÑyZ������DU�^�Q���)�Mԋ\un��o>�d�Ol��D��&�]��_�g��m �$U�oArR�hr�$�<�M(���D���'��\��͉S�j12�Bߪ	T@���?1�T��M�R�.)v@��
��\�H���o����4�?9��?q��}R�'��̯I�����
%��I2MU�� �7�O�?���72v`i{Ձ���p���͍�h&�(8۴�?���?Q�e�yd�'���'���C8Ĕ�� H�1�8A��5�O�D�d�d�Of���O�՚�cپ@�`��$ z�����O��$vN�-�''�	����'&�Έ�n/6�p�*F�.jZ�9���4��ɶP�V��?����?�����B�J�z�R�]1��(#.�rEn�6��n}RV�X��UyB�'0r�'�n�Z��
���f%�OϘ������y��'Tb�'Sr�'��`4b�k��mg�I�R�@k�ʕؑ,5���FyB�'[��Ɵ �Iџ��Ѥr�x�aVl6��ȃdF
s��M��O�cy2�'d��'��I .d+���wdhY�H!O�xYC�+��d�O2��?��?�á�<��OZ9 � A6�܁i"ӮX��'D�'S�I�U[����$�OR���3r����.\�}�jx@�X��?����?��,��<!/���u>1�"��"Ș�+ݬ
jh���OZ�4?�,���i�R�'M�Oo4�VDe�Fe^�yP8�"�34�b�)���?��t�����?�.O�b>A#E� !Px������Jc�0�Ҍ�O!ؗ���Iҟ����?�O�����7n��!0VO޶~�QR�Ӯ�?����<I>�����'�v8�+Dj ��p"�	u�H��g��$�OL��R K����'j�����+�����(U⢑p¡�;	������'(d{3����'@��'�4���'����5��oF�X�+��'R��5 ����O"��ydP�#y�(sOU$�%2�o�*���*s�d�O~���O*�$�O�˓?�&dH4���b"�c�L�q/������8���ayb�'b�៌����Ɖ	�N�8�G8E�2!9�(A2[qh��ȟ��	ɟ�IHy�O_�I��'uꄈ��%?�~��L
 �q(��'%R�'�"�|B�'��)E�\�H�T.Bl��
�睊@�� ��Vyb�'f�'Y��0!*�	L|�É�{�Q�I^"f���i�?����䓕?Ɋ���2�B��&Bō&�@��,�	�'qrZ��z2���'�?��'F����(9?r�͙4�YÚ��I>���?1'@�p�';�� \���c�8.�DyS@)��+��˴�'<�I!W��y�4��I�O���cyª8�H�;���Xg�����V��?���?a�n�'�1��]��إ�LtZp셳�$l�V�Y�i^�J�HF��fH���#d��$��tT:�	�0�t���Z�k@eS^ʍ�돭-������쟀������ݴ&6��'j��O��OT&����(��J�7%�����'D��S$' ���b���yc�<`�B�<W:=���ob�O�L�挌	Ba��(��0�8�
�'�D�27��+t$0�D/*&�@;�4n�"Y�Nħ[���#�W`V�ł5���[�|�I�9Dm ��'�]!F���!��"�^4*Cb�<b�9���<.�l�!oK�X�8��F�|}�yB��m���H�L�hz��ЖoX��Rcc�9E�@�F0hu�P�"��]�^���g��"� ���81V+Z#s�P<��!����	۟tnZ�_�n���W^��J�N-�V�6*[�60X�V�3��ˢI�?	�|�G<O6E�D`�ee@���հNhR��.}j�`Uݱ���҇��+o�6��G@�	S�O���ݰ&`�]zBM��iV�}��,	�%1��O��$<?�њ~��}2�OOk���@�R�fغ%���5�yb��z5^��n҆P�x=R�-���'C�"=�O����	�&��	G�47Xq�e��\J�ĉ�t�R�t��Oj���O��$GϺk���?�]�de�t`�� �T^��gm��+4 6��4�H��c��pɆ�I m������
?l�x�
RBT�{:�7-������v�s ���O$�ɲ!
NZ$ГȖ�*��7I$8~��'�ў &���A�ǭB�����_�]�N��� 7D���S�}v��ń!+��M0�3ʓ\���xy� Y�&� �I*Q�n����RH�2VA	�qP,�r���?��{l�ԓ��?)�O�1�4�D5N6l�ۗo=p>�����G�0<���D	p�hurD�'����#I�G�(U[WaN�[���i��?�Ќ����=@Q˦�'�֌����?Y�4]H6p�,�&4ph<a�#�ǖ8FyB�'e���!%ρ1_E���B�%m�Q�'@�8p�6m��i[��H�+��PjC�[w}r\��� �����d�O�ʧw�
8ĸ4��9W/Y�pu�Ir Gͳ�?����?�Wb��3��� �8�[� ���'�uW"�&�: *��'Y�)9fM���'P���F#� ��.U�H�q�8\�pMN�v��<ccJ�0�x���0LR�'ב>a�/��2�GI_�g\�0�����xb�B�:e�j����d<%	���p=�v�Dԥ�2�pR��?Q#|�+S'9(D}�1���M����?��SҮ�����	�nڞ]B�1!vF�,�p�P��ʹEi�,̓�'*<�E��1'�xҧ�cw��WG�09Q��	��Y���΢uT&q��JI6.ޝ��C	�?!���D��q>��w��� ��M"1�R0ɱH������O�O�����{�N13f�T��e	����9 qOL�Ezʟ 6M?�hЃ��M)�)Y'-A�!�Ԭ��!N�����ҟ��	��ɩ�u�'���JU�%��j]��d}#�kA�n�b<m�)����dI�z%ܥ�&��x�8�ԯ�+o5�&K����?Iu��)q��պ�bC<<��`�%S˦i%��OT���\	�dP���)D�uj �ΉG!��<�A��E�m6�*�Kî)Q�a�}��J %FZ7��̓ѯR�h�<�FbD�vM��1Ro�������$�V��ݟt���|:��I۟��'��$�f��L�f,�C�R��|���fp�'�hs�Q��R��2��+��:lOD��'����2'쑫&��0�Q�$�@�V�C䉀zuLЋ��6~��a��߱}B�I�Z��A�Q���i07�Z./,dP����e-��m�ʟH��j��BT(c6]ʓ	�#(Д2R�
�J���3F�'���'� ���TsvQ�PO�:,��K�i�~�Xws.�r2
�ez\t2�,�P��`p�}%
~�q�S���0@Z}Pҋ���V����3���k��,yҞ��>)K��Lc�4�?Q����'p�ƔQĉʧ�R,��-���'��'&��'�����r�:,E(��d�No���i�<\O�$�=��o�Q��|c�Ŝ{D%�iE�K@Y+��n����O��4��9�n�O*�D�O�7�˗�<̊`�D�/��d��Pd���l̓sl��	�]�EQ�yv�\b-�6�rp���D�U���D��hx�q��.b��s��M	E;�A�	E̓F?�>�X\��FύA#�|�E ��{4n���K��$�P*	�q]D!�u��8��=A��)�)Q�|��}�A��r4�<���H7bu�	;�����L	៸�I��@���u��'��;d4ި@aKǠ$=�(�Z{���o#G�E��	�d��U`�D��0��S�,��7m�(=M���$��r��їL��Ve~�8��4қfn�<�?q����?I���S�? 0	X�n�?S��@�Eپv�F���"Ox����V� Q�e�]d��kP�����<����V�i;^��4�ٶx����c�[�ܩ �C�O��D�OƤq���O ��s>�����O��G�����,sQ�8�c��uݮi�퉄P�O�Q��Z�m,��*"!@����'B,Ă����$W,->�d`���,-8�K�N�#�!��L�Sw��c� �1�`��͒8ih!��
�>x��ThƩV�lX����C����}�Q�	�7��O8���|:�)Pn�M����e�"��ӎٵkbU����?Y��3�@�E�i�1O��O��95���Q�*��G�5Ūl�Q��L*z����h���< �B�+�-�&^\���䗗%�"�'��O �SM�$P񎑼�8��@Jl��A������<*a�"�!�@m�~���$@x�M�D9�+ƧI���W刄Z�5�DA�v�`6M�O����O󉓁3/����O��$vӤt��G�<�Z�P'�_�[#t�6�Gޟ$�<��ҟў���1���TK$2x�RI���O�E��O�Yq�R(e��yPE���+�8m��@�ԟ��<���>fA�'�E�戲\�Y�F��V�<A�j��L8��jRLբ�����}�.�����M��&�(t���Uė�Tp���˘ҟp� �1�|y��ԟ��	��Yw"����dG�D�P�C��Q���H�EϾzv$@���% �4� wΒ�t6T������ e`�@�� ��l`ph�8�舊��ȒC�^�1Sm�0��� �"�Nڶ���e�{�F̂uM<`%n�~��'Fў%��8�	Ă�� wAO�ILg./D�`��l��E�!`̠�BA��:�Q��S�Oh�?���R��iޛv*C�+er��[bL�
R�@�����O��DT��6��O�瓊U ��D�>�.�:ZR|��a�vf� �P^؞��H �dZ.�]�F�E���x�p@��kKa{����?��O���MX7P� 1&���%��"O�DP��CrDt#gD��@!�lq`"O(4��MW0m��T1��ή(�PUB������'����yӄ���O��'Q�T��D�S�a���ee(Xg
c�e��?q���?	E��++f��7�xZ>I��|:m�v(�&D�n<���R�WY���>����:���Bڼ����~��.��n�2I�g!_�+��a@���a�g�1�����ܴ�?�M|R�d	$e�j�ۃ��Z"`U(Ve�uQ�	Oy����剃9�0�;���Q.�Ĩ� hd ��$z�Jn�t}"bK�=hā�C���F�	PkG"v�R�e\��E��ٟ�i>	��*ԟ���֟,mZ<8Pd!�)O����c�jt����'��3�%O��f䎏 ��[�O2L|z1�ቾ�H��I�pp�,����]��pnؑ?�4�*����'�<"}�':H�ak��B'f�V�V8E��'��ӕ!V;M!|�ZD}{B,S�{RA"�S�%\�,X�KC1 `�E;��q�X��=�*� `F��?����?Q�!a������	�Z���r�[�1a�E�I"p �f�-.82�`B{���;�ޠ���(�Q�5��!�gӸqb���9�n�	ߓ�v�!6��3&�0n���7NW"��'Z��'����%�R�
��L�Hm���y���sE#D����� ',�[(4@���@�L&ʓb1�	Oyb��`6�~��( S$�����D�	!�!���џ8�I��� �����0���|�W�џ�'a�Q��X%a4�����Y���=Y�E\�I�%�vT$k�)(�sg�8������u��P� ��GM�5��A�E+@
`B���/D����)
:o܌k��!�^j&e"D�Xpf�8A�q#W"
�&��P�Ch�z��Oh��F�^�%���p�O�^��"eI��\��gG�?/<��P�/Y��'�#��>��T>�Ĉ& ����&Ĝq�*B��Z/5�O�����)�	�./��M����8dX�#Ċ`>�O6���'��?�qԊY,_[blh�%�/4��A��;D��!�!ƋQX�=��� � 4;�$:\O��=��
_7q��X0�dH>dҘ��	�;�N�1�oӎ���O��4��)qg��O����O|7�C%xiH����]?�rWK�)0�����O̓���A*��5��,
��g(߻UNPy��$�q���� �QlP��eũa`�h&�)�
 �	g̓*��>��n���Tqs�}"���-_�t���S�? d��$C��0�4ؚ�.�6������h���+SI�ag�3A��u
�D�%\�չ�'�����\�@F��'3"�'��םҟ����dQ���1m��)����q����� �sy�����:m�������Zuh"�f�M%�6m��4��W� t� 0�6�'�6��)��?��9`��?z(�"o�*�4���O��oZ�l�'�B�xҧ]x�6�RKW|� ��s�%�~��'^����4�<�C¢,=�]�0��O��OZ��O]�<j���(�4�M�WD�j��X�rlS2O48js�Ƕ}vB�'�򦅝6L��'���T�T��A��<��R0(G�8�@8lO\aE�xAU��R� Ղ�=��`c�K��=�G#�ޟ��'��1Ò�͵^��R��Ԟ�
���'�!�OT+YHp!��ں+&ec�'�z@P6��b�0�c�*sn��WI�{�f׋�0�M;��?�(��a��`�<PY�%X�-� &<L��Xc	p�D�O����YH�$7�|�ɗ(�2�Q�;`�B�`r	�5J^Vc�@{�>�S�S�Aϰ��oΜy�X� ш::c�`4��O#2.�sd����ĀTM�P����`�<�RI�-���#2Fٴm+�`r'�R��p��{��\�[��qB�!V�i��1��!(�q�l^���I�x�i>�����I���o� #�b����\.}|9��l�;��!���'x:�3ړL��(�1o�7h�^2qb�
*�5b�ቲ�H���)G�$��#h�Ui�ef�P���b��?����?1�(�g}�j�6CB��/qqd��%��$#�O6\sQIʐo~�#�3x;� �d�C���	j�v���ԯD��{��(T���Z�oGן䨡H�Z�^��I����Iʟ�s]w������P(0�}Z��ԝ6�p�3N�4
4�;�_�5"�]���e��ܲrҡ2Dj䃢M˸&~*X�A@x�j�g���Op|̀�⃙��<a�׸i���ơK#y-�ա�B��
7��O2��%�$�O4�D%��̇/?\�G�L���q��kI�g�0#<Y�/�gyRC	�U+�D�K����@��~�A�6��$�b}]>M�g�>�M#�421L�6DF�n���{(J#3~<!��'o��'��2��'�0�R�'9�Ɍfi�I:�'��5A����:I"��D�8>��'������-湸f�X($�&hۓ�L�IG}B�7m�~7�S�Tk�p3g��yR�"l�d+���T�`������y"+?�*́�!L�uꠦ��-��=�>�C&rΛ��'7�Y>�g(�� $��Lt}��{�/�9N�]��ПD�	>���b�U�S�����2�4�d����@�0!F��>��A�QQ�*��U�%���BehMQ�޼�g�H�4���I\�OO�q3�M��-ے��v�M��'��1A�D�\�d!B�ק!�V`pד&wqOj�I��D8w�����ʋOMX�h��VYݐ�{ߴ�?���?ͧ`��t���?)��M�a��M�lm�����q"�x�.�&+���H}F{��^�)Wh���'��� �ٻ45 #<Ae�>IEMX� �6X��ߗ!# �	rC�T���i����\87Q��b�i�i��
�Ff�!�d�,Y��lz���:W����E��qO� DzJ~�eoV�xv�3�+Q�^�����Cz�<�ʀ�s��H��- t�0���r�<q&צi�@C�ٯ�؝�ֺolQ���8���"��rJ�0st��a��q�ȓva�9��aց\��Y(�a8HL"T��US$ ��k��t@���g
F�ȓJ"�I�5�Ҷ
f�`�e����� ���X�%ִN&�X2/��d�@ć�?,�e�&*�0"��BӘ��ȓr�q�Ԫg��5��H�K+ԁ�ʓ2�8=��F�vp�m�k��y�DC�I.�����I��>��@�Q��B䉢2=�����݈��1�R�&ĦB�	�K�uI&h�7EDIGc��G�TC�	% "Py!�C'*$�a�Auw��D4 ����+�x��t��?o�!���*ab9R��]H���3Uy!�� �9��:blV��S�W�V�#�"O��˳.�^�vqj���A�a��"On�ٔ@�%#��eP��'wF��xw"OVH��B�5J�
�i��<�.��"O�����>w,����5i+(���"Op�ҥ�]..m�T��+Z	�aX�"O�3�ń4^c.=����։ؠ"OT��fQ�s�"8�/[�X�x	$"O.�9�Kp�d�hP$؜7��X��"OH�a�'��K4�(�v-��U@�"O�H���f�ЄB�k��x���"O*-�#-P򎵻�e���a("O�u"gk�
����J�n٢"O�G<`�X9rD�����"O4���@�&hq���5��0H��!"OJ�
�'�Q/�0�mK֍0�"O>ѩ$㑀=�j�S�3-M��"O>�2�	Y�3�L��5�/� �"Ones�oR�0��oܺn|�i��"O[�_(y�����Z�c��e)v"O�Iˁ��1).y�EP27w��f"O<h kʈ�v�1c��[�݀q"OL�A0K� `����-��Q��"O,H5c���|TI�N�.Pu\��c"O�p��@�0�����oV~��+"Ofx��*�7�ĘX�d��TϦ�8"O�H�F��-7� Z#�37�"�$"O �b���k��|hT��>�y� "O�0`��Y�SJ�"�h�;Ӥp#�"Or����
�_~A�Hn��}!u"O"j��O�c'��8��0�j���"OH%���/^��hB#Z�&���c�'@L-Д�L�U��$��7V�@��!�'}B���ē��|�'��/fw��5���yTLF~b�Ӽ;�v!������b5���S�1�ÆF1@�!�dX�<��Ie�C:M�pK��޹a��d��i�u�D ۲��)�'}7����01<t�R`����ąȓO�d)(R�W`I"�k���j�O�Т�@V>���� �|���!V98&���#4T���� ���&ײ����c� � �先�/f1#O��#5��k���5m�oN��3��I�Pt��F�*^�1��U�&��qt~`�ˋ�Q".�i�"O��QE� �*��1A�ܩ 2@3�O|A�Q�@1H��}�ӫJ7Z�>�ȥ��=V<�;Ј�^�<��J�##3����[�SI����e�\����� !E˱�0<y ����a�`֠���� \X��8G&����!+ �ΨB7� �,p*f������܌����Ao_y"�q�+G:��Odl�EUx���>]���R�uX���ۛq�����(D� ���
��u,W�*3�a�'Ϣ<QTV�]��➢|2Y���7o�}��	0�D�b�� �ȓv dR��T��K�� �ZL��C�)�D@G"M�Zd�0>�LфȓF��]k#=4>��
���U�&����p$S����E�⁗�99�$��D��/rqO��8s�-RP��J5:��P"O�(r�aC�(�3��5h� �®�b��4l�4ڂ��|�j�;a��t�����" A��x�*�:b*�p��M	�
Gh��W� x��ɦ(ؐD��I�F�̈b�pR��C�+�M����$F-{̭�R�#��ɽ;�> c��._��+B�X�;QB�	o���e���~��V�? ���	(z�w-��|@ӧ��	����h����
g���"O�TӶ-�KD(�[Ui�2)H5�4��I�J0p,*P*-�3�)� :�z��U��Τ����<+"�i�O>�B3%��g�aP��ܫnR*L���U�'�*�f�PT�ʵ��"|O�Lf�Ȟ'��A��K�~��s�'D�$Y�LC� ^��� l�2BT�6�3>�����B1�uQҀPi�!��>@�v]@��<J?z��4�Z� ���)y�r�8�Ҵm}�w���
)Q>��g�͗z�J4 �j�
t h�l D��УF��5�d�Apd|�k��_<;��04I�2O�Όp����}&�`R���Q�4i #ڋS�~��a*9$��:�b��mK����#
�g(l��J�6!,b`ʖ�ʺH2�`+�b�`����D��+V�4�1�ˢx1���ũ;�Oѳ�F-H�py2WNW 5��%�4S�~q�M[�A�!�$dl�a���G�}>^�rT��p����7�x����=�H�"C�L��Q>����ٲy�rԒ'��.�	� &D����
Ot���@�� 2
ح���Y�����^	&b� � ��J{���qO�3�P;b}2,A���g���Z�'*�D��v��Kc*��
0�B��r��P�^�5��p�] eo�z�f�"��qk`K��'��@�!	��O����^Rp,�e� ��B@q���μ��#�8y�#
���"O����ȗ-|8H5�� �9��ET���1���ڵh��X.#�Bdr��Ӛ#��P��
�#\r��R�e�C֖B�I�$�9��L�I�Z��L�]}��O� �E��V��t%>c��@FU�+\�<q��vގ��l&�O���)yȄ���Sd�iP�Î�b �'�X ��?7�#���?� �Д!�U�'<	��OL2;� �&H����$�ȘX4�_���$];� 1a�+D����_�g�kń@�T����`�>�Ghت%ļdN�&V���8�'R`~݋V"
x�(�cЀ�q3�4�ȓ6���3dD��c��}�֬� u�r�x#ș�@AH�+̝7k� znGI�3�ɺO������L������L#]{C���N�Ѐ���*�&���m�}�h� g��)��	��-�|���ۓ})l��S��t#�$��%2��ɂJ��aB�`M+���Z/^H읻A([1!$i3�Q<�y� R;X����'�=K�씀��ɩ��'r^$i��@�s�x�E��Λ�{�D`M�ΔȦE�y2a�y��\�r�΅�0	���̧���wL7-���'�>���&�ݘ�&1�>�Aa�*H>B�ɑ$�q�CaѤ
V���t��	$hb�h����:]��E]�K2�P
ۓFS�@3΁�j��$P4lH� �F�C͹O�q� ��"NL�P�Ժ#�ʜ�:�����E�2u����Eq�<��
ӸA�X<���Ӄ�J�(FeDF}Ң�?}� pj1+'8PI�)�`�O���*�pP���H��
�����'�N�(Y�En̩ƭY�My�h���ġ|���Qܴ8Ѵ�i�NV���'M�r�K,q �S��Fu�b��� �:\fq�K�J�D
'e~xi���%��듈�=������Ft����P/7"䡂�mգ=�y�N��~2Om���0���ZS�?�B!�s��4KP)r�}����2n��q�E�1�y�	5�B�Q��M [w�5��k����D̃Gd��s���\i~�ӺC� ,8���-O�:%.C6=g��J���&��I3�'����"�Q+u�h�C#oE7\Q�9G�*tAwyyb��-D��갅]a�'���8��I:��30��30��虋��S ic�8��dOLJX (�ꛃ�>�27��|\УPN'!��1 ��fnT����-�h�����>3�(�H.Vt��	�8:�J�j�^��������O�����uf�;�/�$ކ8��'�
1:W�Y@BB�(I� ��O:�
V<�,H�p 5H\��k�v<If�k?���< [�܆���/V~u��7%=�p���W�;�D���+ޒ$�Tas�
O�ţ�H;$��2�ǁ�-�x�0�D��4��7/
:!Ꞙ2p�8�ӔvT�3&2=���s�d��UNnC䉦Z�Ԑ2��J��p9�[�$v}��ɍ��h�����?AB�7�gy���<7pl�F���D@�!��yR�9>���C��E�b%&���b����c�	8g�x�Anֲa#�y��M&dŠ�[��1;5v�*w%��0=a�K��1L��R��>	�
8#��i
��L�șQ���1��'�Ƞ����>Y�; �Td�uZ�V�,)H in̓W�"(��,f�I�
Ҷ��tY>%b� z���=��U���ɿ� ��*�me�+��=;}�W#�pja���ӶT=�CCP{0�Yߴ;2h��"��Dc�sd}�����UΓ{�ܤ��H�"HR�0�c޲
����ȓ�&Hh�B�|P����k��/=�!s�/�0!���wE�
�@���CX��(`�'U���K;-;�=ϓ���y���HݓD��� ���	��a�!I�]\���/�<R�>�2E)�_��,m�ʄ����*D�R��T�a��8��M�M��jT�I�*�xAS�T�;��=���D^c�8����CRA��(W5bF	��ސ_+Z�ͧ+�vm��,-� ���cӒ	�d��JS�J���jN �O H��O�]�"���B��0�#Ũ�jm�����"�롈B?P�$�_�6�����>�0�;�8 ���)'a0����Il\x�"Or�X�JhǤD(�I�Q��3C�F�'h�<��LˆT�j����<7
p�@Ҧj�dhe��T��S�0OĥXf��V쀀�T��-��E�T�'B�\��[��u��E�i��iy�@�$�Je:��
�g�|���˙r��i;O�xRf/׍}��A)��$C3�8'*�f����M>��'g���e
M��$�hCl�p��H&JX����f��}���S�`!2���^�I��$ڶ
�&j\<����j��(����G	HA2��ӱ:��Y��苡�3@T%1�6����|���S�� �D,�.�yҗ'�Q��*�5H-�lRdBޛ��x�D@5_TؘH�ˑ"l��LH�n� �L�5�a���	J� �h +@�ݨO������e�YA���<�R-���'�Ii�ƒ,9�N�Dk
2_x̉��ʑ)p���o[�A����*�)�!�D�\�b�!�o
y��TSH @��'��D9#H��E�~�M�6�|�����6>��,���Gw�ؑ" ��'�!�d��H�(�@m�� ���ʴ�+L�fl����I�*Z)M8��T�I#?����/KNɠFjA&r��Ћ2nh<��Ŋ�f�@��J�E�<T�g �W^��[6Ń;��	�ʂ�yÓk��a�� 7Y��p���;qh���	,PN2E@�c	�=��`��'M���B�oH�>�R��,]t`�
ORe��FLx,�lD�y n`���D�x$dx�d#T$YxzxJ��G2ܸOB09���	wE�]���M�|]	�'j21س�I1G��I��I�� ᆓ�>��x!d�����(���5#�n0� EY�\q���4#�P<@B䉎!�`|��JD��`�dhʬC�R��m\�N@����!J���2˓K_b��6�J�mf�`w
~��y��	��H�b���1���21OS�Br�	ԃ�n��3aFE"��D;ռѥ�|ޘ� +��t����@�u�q ����� 	 {�|�BA`��v�XC�I�Q$n`�u�ó"|%��i�27���l�up�{���i&X�� �����o�<Q�$���'N�i�*
%�4�qj�M�����';�@ H7Q�N;�h�+`����'l��hP蘮|KZU�1$n��*�'2�0sʁ>�B�20�[@4��'�P��`~��Y���֋w����'��ۖ��*`[��R��S될r�'��x3��Ϩvt�`qƗ6f^�U@�'3j�٥�M� ��c�^ddڹP�':�I�h��'��a�2��[N�2�'���
�0�B%y""T8z}�%��'�|�%Ȑyc֗�H�Dm`pn�<тo\�U?@yAYJ�T��y6C��1V�d���dO�<Ȱ�rR�6U�B�F��
�F�ԪP[U��c��B�	!h� �Zs��"d��갪��W��B�ɞCS���sO�jkDP�.� \���A�%J[��x1'�À��x��Bl����	'D���'���F��D�C�®bH�R�(D�0*PL�;�܉C&튝^|��''D��(�NI�
%�L�3n��h��e�#D���T(.P"T�I�*b)R�?D�蓶Au�:懦Z��G�1D��9�F��7@G��<y9Ӡ0D�@��/)&�=Z�,D9�29�1D��2����_�f�)Q�Bc=0q�(+D�(PC��6X*�	E�@��>�`��(D�� ^��RQd�9�I�//+^( V"O���B.�a�6���@rl�"O�Ya��((S�r�˖�`M��S"ORI�á�]O�}x��H��R�{�"O^x���"'Vx|a�g�(�z�"O��j�/�p'ja��ա4S���"O���"Y<P����,L:@���"O �1�E�/'�B�q7���N(�"�"O���%�ħF�*5��]*x�K#"O�e�u.��g�f$��B�����"Ol�E�B�.cȝ�⫔��Z���"OVDȆΏ\E��� p�`+2"O
��# X	^B����Ք![����"Opq�KǠA7�#��9<<&�R�"O"�xTK�>���gߩ_2���"O� ��@�;���  ��7"O��@���C��4�&�WAk��`�"O�x��H�){ b��ܻ@LvP$�'`��y��.
$��dA�!�\�;�@3e�� �gd*�u��U�c��~��΃dLB%`�5U'(h�*���'�r㓽�%ad� 
A[��8�S�FS>#�J0ATi6��0��U��y���*����_��5�Ǘ�hk��)�
���P��qaL#U��ɔ��y2C$!IR0��䙂�K�aЄȓ��S�Z�¥i�P�w�8��Q�O��?�%L�6��x���ZE�ň��^j�'��9jub2��m�0��6���#	�2[4�A���ncH����lًG �7�T� ��� ��$Ȇ�8����D�k��@QV��F ��s+stqO�����z:Y���?04 E���)Q�6� �@��p�T����:kI!��5��1��k_4.�4��&k�+��@R��=�D�vG�-,2V��GT�VY��X�Ɯ��E�֪\�Dc!򄓺g��L�B꘸`P�Y�p��"P�8��4n$��	m��O�J( Q���'F���
4+��q� 9��3A.\OD� @�:��M��K 8jlU@����ҐCQ��D3�F%49~l3�?�%�%��z��|��
�u *��=i�ϕ@���U%��X��!����'z���ʡs#V�3d�
�܆�PZ���P�!<}�ق��M�/��� ��ٚO����ύ(X����S�OT���ҴA�mĠd���O�t<��dWF�q�@]�)�H�@�n[�!�B�7��D�ֆ�+$k���H�
d�F�G|r!�7%��h��`�6e���CЬ�p=��E�'7���0�ԥP_���!� N6�����2O�T�兘]�	�`k>�O�������}��*S&_Q$]�g�$��h��1���~�e��ˇʟ$E3'��jD�kSɉ+)H,QV�Ĉ)!X��'��� P�<>X�)����?/`�ѤI�� t�狅��8�����(�`�� A�=Y�d��EPM`�T
&=�Ѐ�WO�Q�b	�Ew �Vo3~�М�'n	�r 8!uf1�# �;b��zd	���S�g:
�'��P�6$I�k�vU��ǌB)���דհ�3g�@*(���F)-;����ɓ{���!�͔|�аW�������Z�l%�"|s�Qs��d�g�@e�$�qe�Zܓ>�9��m�Kz��.C+��)�)� ���>���xfH!�IP���|nX�%IQW�g̓��}��D\��e�pg�?�:�i�Bȧ��`�ѡK&H��@��S�Ob:�+@Jمx�8|��S���sB� ����w���?)$�5H*x��Q�M�y	j1`6���?���G	Y�[���#&�jׇ ^T0���BW#v��O�������a�qV2U��'�j��Q�ܤU����K�}
6����;%}�	;U�t	�`��E����e���:�������S
�C���k^��j��P;]���4�q��wzQz���F0]��O��-Kx�pJw��܌�r�.ՠ��c��2g.Ԣ��x�IҰ<��d��
�a�m�n�{$�w�[�n~��BhȶiF ���	�K���ɶ�.m(��H3�.B�P�3!
�h�B�I�mi6�3��	?d���'�"�����M�� 	Ĥ�}A J��x�����g9Zd+��4H`�y��  r"�|���C�Ȉj��I���(��Ó�o�čв�ގ���T��b<)�,ٻp������V0j����	x�'���)�$ɛ0�����FP�'>K���@��H������7���/����s��6[�$�b���ZK U�� ��}Ll�QD����S��?�  9�s�O�N�~yEJM��qS�"OT�EE]"zvp4�b%g@)�1�Oб����Uc(�9BA��0<is�`�fl�����@Q;�,�M8��A匒0�ڝ��C	2T�q���O�}�[�V�	%G0D�"GO����:���� �q�0+��	�2�����6_���������mT�mw4��p�O.���^������K"o���s@����)C�X(	��%�ۡ��IX�ű��>7�_9�~�ľ8�ĵ��W�f&�a0e���y�혓D��x�˩Sjm�����yҷiϾt;kZ�M`���g	�rM<)feh>U�RC�tgRh��+�o1L��dn2�O��2如�	����Q�$e��3A�X,N|ٺ��,3ORnI��l�-_���Ƀ|��d�	ǔ���풇{�6	�f��}ܖ�<��e5NG����傧;r6�b�����gBR:4L�
m�������@�D��#㟨҂`�8�a|� j�N}cv'
�"����J�� �b��&���*��ڞ@��%S5O^\!�/�>	�Ӽˡ`�6zE;g���Fs��v�<��%I
w�x-2�E����P���8	ݒ�r�'H4� [�H���<	�Ī�%JX���Bl�9)� ;j�jL���Q�
�Pz��)�O*@�I
g��(�3�0ZM���qɖQ��LO��y��'�QZd�?G�5J2�1pZLً�$�;UI����8MC���$���Q��(%%�ɼ���þ��,��VZ��� !��Yp�E�E���҃�2�`��%�ԹR��'w$Ik�b�@ʐkg%ؠ5�5[rG��&�&����6ւ�U�H�e�4h)B�|R��y��_&�@P;2��<rxQ�N�?�y�F?'�<�!)�1'V�Yp�}j����
ϑ��'�r޳_qVh�Eg�lқw<H5��!>g6��	q�[�0~4)�.E��KԬ /�	d�ܪ��p�$�%q�=���l����/�"xP��#.	�`�̪Z��#<�qf�p�YbG�Dt�vIu�'tP�un�]�p�[fO�D�t�*O�d�Q�?5�,����=@��t
��]6\��Q��+nAa|/�Co����8/�$�5���`��L2��P�܀�f�X�S��d�O�n�N���ZD� �p�,G����u"O4��r��x���-nðAS� �h��d��%;��5
�isލ�QN
O#NB�P� 9���'&�O����ʗ�Xcv��Ǎu	�sț�.6�Hs�Ύ8�y��1g ���f+�gk쉱��#�uG�:H����#���i��}YVcm���<��E�F���'艷)��dny"N_�5�p�S&�<^�0UI�Ɔ�'b��X�4
xڄ�G�'8��$�ɬAAє�5a�|�[��*	B��i4ɌQ��e�1O�pS���!0!7�v|���^�Z#���M��y�j��u�^i�����2)����?Y��D�Q�Č#�B�lL�ړAٿ0]̻1~������j���)Cx�}�`�~~�hё������=�1���?p�v��C� �F�;�A�WI�i�Ǵi�UA��Ī1�>��"�-r�����^��?!7�΋C��9��+G��%��2��:@�OX8(�&�u����S�ڰ�)�TMC�"<�)С��g��j%�4SU4%;$�S���8&�'&����j w*�.�aW�k�NOǦ�O1�B���� ��̥Az"�[`�"���V��`u��?��f��7���$
Jf����iq�����P�����[��z�Kp'�O���=��c���� ^]�<��CM�{�n¯#����녁uI��	ʱF�I�W��$Ӈ.  hG\����0=��g����PL�&'�7*��U���"c��m�m��ĳ�
�j� �Z kܑ}�����'/��OR�����mEK]�xju��HA�`��A�4U4�����&}�I��-"h��~b�@BEf���&Ζly�{��7&�$uR`N_;n��L���y��/	�J��6@�$'(�0E�H�2��@�Id�'��y�P?��!����!�+��2F�[v�7;1џx3����z��fəb\�������A�TW,[�x�B�-��"2�}�I���'X>�S=,0l,�U��8>���'b�˥
�Z��Q� ��k(Oj0�Ba��`�Pu2P���Xvb���Ϙ���š%�R ��%�=E�!�#W4�ZX6$"i���Q@  2a�rDqt�5�Hx���ӇJ�X����ʅl�������J�0|�ԋ;��'j�$?5������������(8�^�)%¾�x	�!����%X�f]��P��_�lTB���b�E̓,�B��H�P)%������K��)1c������i"^�g �p<�gL\*��z1�A��'B��p3U.ȩv4-��ݴ14�y�O�I��-�hM�D �3.&�;�ʞ�%b�*O�-������b)b|8)��>"�D�)rV&ՑE�����(O^��L^ɣM=}.L���L�(09*�앰|Zd�����?(	Єɢ����O8�3ei\"}��(���>��]�u���$�sFΩxP��Ĕ�gqƄ�5n])sL�#g@ �i�,�:�gM��p?Y���L��Y�fT=3mN����#N�ay�.݈:�ڝW%�􃐡�>��b"�z5�I��)�l��Č�.����6ƖQd� ��ۂQ(8ᚩ*dїKV����xR��o���Z�-O<�P!/L��'�lY��T�p����,3�|s��m��/���(� ΓM("u�dC�7��	�]��t���� ; t(�� }դ��aGX�-�~��P�"a�zrυ*T- ċƭ1��,�S�ޠZ��]�vI�" <h�7�"z����	#}�H- ��ȟz���'�ٻU&fB�Ɍ�$Vm�K��M���@�J��EiV"@�����' (P�&3s J��;>�n���/٦ly�尐,K+c�>Ї�ɅOt�Źᣖ2���rJ�S�6u���G�Nd�d�s�М�4�,��u WC9.�FQ:#ݙ[:��ѫ�>yԏ�
C�&l(bN�6s�}���_�'}H�2�gҦR��k5��7Y���z҃��6�Eـ�X�4p5�ģ��[� �)��I�M����EG�
�
��%��v���>�@�ߑ��KԀ�.N�B�Z �Er?���M�F|vp8"�2Q�H#��н	8\ʓ�ĽJ"���c5
��U"W o`ܤ�%��"mpԣ�,Y-b%���8���0e�2A���;��
+Ae�,���֟i��,�B��?V��"x����4m�0E8��y��!�:� ~]R�"Qɋ A¬�T��+| ��:�BX���_/\�,�!�/�<Q�ʅ*���7Y~|�ç��"���PáE�6
Y���G<z��"�#�1J�)����M�$&Q( �E�7F8n&5�k�b�'!$�ꒅ�*i�b���,�9J��J��_"�}A2(Ƒy`�Ͱ4�G�iwͲ�j�5`b�N�,kj�����.?��|C���8-����`+��n�݃�.�6h前D�`1���,�X�'BS����	f�w`��p�:Pb�uh������h���l�����2@�h�	�������7H���h�8`a`�ІBA�}0&���+K� 
�-%8$� �C�H��0`�:di`�ԎR }��n�'\�亗 �oBf9��8|j���,HA�����Z�A��V�ӷ2�ܩ���]�.��D��E��\h�bӯ^A����B�!�t�P�ˇR'&ݪ���S> ��eWr���J����דD8D�gؕWòL����6���{��[|F�0�a�(Q�*�U�z���o�(��R%!�VW@�y剠9�ȹ�cٌv!>��̆�_|��K`�̟i���:�L֥}�����3�c�/�u`T5$2Q5��:9�h*1��3%Vu 'T����	�2���'	��Lb�MI��{0��)��P��"jä�J�DO�2y��?��w�qJp�¡_��$��%��d �'cr���^x�=��d0�5�'�|��SN?s��Lb��6`}x�'�zh:��UР���)Tˠa�'�reˣ�7@ڶ� $��K�t��
�'BH��&H��2#b�:R~���'n&슶�ѽh���r��z5��'T\`�E�BBP�!�U�nX�Q��'�@,�����y]vR�ɲnCl�c	�'�<% ���9U| �óf8�iP	�'�@}��(�X�	�j�S��+	�'�]��q24!3��J������'u����_�HT���2�4`�B�	!F$�1�� P�u�X�wo�$��C�i��U��d��v���s��C�I��p0�pF�4S�l��p`>wUxC�	!=rP�p�k6&��*X�WjC�	�28\tZd�����3�d XC䉲l�R����(Sq�Q�?�:C�ɠv>(�.��K�� yCK5O�BC��%G��`���Źd� 'ĝ�7�C�IG���u���B�eY!N�B䉔=o��b4�ٵP(rD;��U�Jj�B䉵f֎�CR�_ �
���U��B�<1����b��ӈTВi��dZ�C��;��4H��3w�~  R�3py�B�	�J���Aԣ
[0T0s�N=�vB䉆>��]{\������l�ް�0�$D���-C�d@l�+!�ϋ`�$�2d#D�t���%���JQ)�5h(����?D��#P�>Hph'H��o�A�#D��W�O K�����s"�t��#D�dwj�(au���Z16��#�"D�`jFP6fV�����]�dD!@ ;D����U�߆��f��k�H�@N-D���a�^=H�U���+hJ؂�)(D�� ����7�x�C,�;LX@�)D�� ܵ��:QP�J�d���9�`"O��	U%�!gPA8C�
+�6��""O(d����ӽ=%�eE�8�y⠆oπ��0ύ�A�L�%���y��M�N�^H��V�h�@��Ҷ�yB�ǝam�h &x�x�g�
�y;����U -rn�re��yR���bgFi2kF4���9��H��yr��&*5�S�>��)����y�)�P8&Qj�����t��1�Z�<���U�cԸ��an^�pb�0��DM�<I�C/j�D�0�C�##����BI�<"&�Gz)���օ(�ܩ�`�H�<9��k'b̓�� ?<�(-�D�<qu�L�_0�A��k�\J��H ��T�<Q!���Z�:��N3D��3���Z�<I��L�Of$��Fd��E���C�L�q�<IQ(H=W9�UYD��(HN�V��l�<IL�9pnĭ�Eb]�A�@Bc�<��E��|�h(����WJ �4��S�<y�Վ,���u��:yRV�����W�<��+^�%\��˲(\�3���`f+P�<I��בDb5q�@�!̙��7T���%m�a�I����W�=D�,�cnOt�
��!-3�,�3E?D�$i@ff��	Sn"L�v��b)D�0��� c��l�"JT�Hi��<D���D@�>Vt!���="tD(v�8D�lP'�\�Mc�,ʕ%��������#D���G��%�f�bB�E�c�t{ǡ!D��0lC�> :0�ւϰ �Q��<D�hxG�1sO�����)����'D�H�.U���#�N�.�j�3 *O(	C�k�m�(���ǽh��2"Oā��EQ��p2�X�(�jݩ�"OVE�+2�����L����"OJX+�B_
2#N����O'�a(�"OL��kX$��#kZ@����"O�t�!�W1�"�+cI�;%���"O�i���G&���W�Dxʱq�"O �;F���v
�1�&��?EZ��'�2�"�( F�0�Q���'��m	�'�DI,�d�^�iQ.��)�����'�t9�@�"<#�D�0��"(n��'˪����+0�8��wK����y�'I�3�j��c�r��'%�+;x�pB�'�-��&A�<�t�A�}8� �'( �rg��*ato %dP��'�2����8B�{@�$(���'^��fð;�ܹ�DAB�m��:�'�8�I�V�Z�6P7�_�!H�'L
)�
A�2}��¶Ok�<h�'ʺ����=bT�� �O�:�'� ���EL�1�<)�@
yKA��'*�`�Q���q`��ǳu�@�'���!��[6@�R���j� D�'/�a��%m6@� �KhQ�X�
�'���@B���w��	�ℐ7ep�I��'3�kP�$�*+R'��*��`�	�'ߌ��qJٔ8��
RN��VzJ��'����8Ͳ����2���S�'<t�4+O Y%���eS�w(�a��'��D�ʂ6]8` ��ț�l�PB�'�!�P�����=Ӡd.`C�Yj��� p��7:�$SKa�H컔"O��B
4H�~�
s
Qk��0"O>ŃiQ/[E�@;��>��т"O|�����8M�\���D���T(d"O����4&t�Q c���
$"O&�!GR#�|���KA�ԣE"O,1ĤZPB �B��\C q�"Of��4�M�M��!�5a��Tk"O��,Qr�q�ɓ	D�TaAD"O�C�E��L[`�s�ɰ4I0Ԉ�"O.� �LѾ(nZ�q���`P�!�"O(- �M�p8�T��[�cD2M��"O����b�@�0`A�N-]S~U�g"O8mY�<N)K�	'?I��"O6���+�C������
"3d-�G"O����ζ4`�=�墔�;!H��F"OBi('�Oi�<C��42�ԉ��"O �	�ؑLF�(��D�`�>��"O)�����L�*�
�2��s"O�)j�X�V<E P�M��J���"O0�xR(��86q3�^�'���"O��ہ��1aPn�SҮ��9�BHe"O�1 ��"�p�H�q�"`9�"O>�uL�T�F��VN Y���v"O���0MD�k���S�+�C�&�1g"O�)�C�O1?���Qjë]�<��"OЁyb#N���u�@�l�ꀒ�"O"�QF*I?$ΰDcu�(dk����"O���@���Bh���.P�����"O���C�;@�5�$�ǧz�B�x�"O�T�o z5���_k{���u"O���ㄫ��0J�'��KFi��"O����[W�8�Bf��n�V؋'"O`}C&�Y�/��arW�L�QaZ�C�"O�(�%��	�,X���>d��"OJ�!v�!͂]����c�`]i5"O
�����,@������̋:�A�g"O��ZPA*J�мq!��:�"�90"O�h0�Ћ>~\�6��k�dr�"O*��S��H��pp��W�v��"OZ�`�C�f���`��o��x�"OH����,Fe�`�L�u�fU��"O��*���0��D�s���3�"O"�{2�Z�s�:�q�ǟg�ŉ�"O���eNЯ_=>H 4�Z�0f����"O��n�-��tz���/FNC "OD�1g�<S�jL�\%3�A��"O2(��+F~�3@�Ű�2��"O Pp␑Ct���6!� l�|�D"O�(��%��e�fX���QJO�`g"O�M�e/W�(��%�v��8+��2�"O�i1䙇\=$��4Md�Qs"O�IC�\)�2�X�����B#"O��ۦ)P,Q���(c�J�e�ME"O�`���O��`%�רMCԂ�"O` 
fmY�
zm��`�&C`<Y�"O�#�3���`�]����"O�i��uɑF�Oo��a�"O�=�6'؍��)S0���y�8s�"OX1;%J� ���Z��yHx��"O�����\W�M� G�
��"O�!�Ԅ�!A���n°*����"O������H�5)rM��4C�"O�E��*�$z?Ҕb �	��L�z�"O� ��KQ���Hs��wM�W��%Y�"OV9�@�Χʚ���^4Du*��"Of�����<R/�ia�'L>.h���4"O�l�U&��i�>�q�Gɋk�� �"O8��C��#|���4�:��50D"Oba�Q!E���
�%ܠ%l�"O *���8&bE��Q���2"O
�
wo+�����c&M���	b"O6̡d�O:
I����K+d��Ia"O쉃��ʡ���k���=�>ɐ"Or��s�:�����͔�!����"OʔK�n$F|aس`�aH�"O\l�a��+��<[!��-%��u{s"O���q�"L��`W�L�N�x�"O*��#��_F&n�W��4J"O�I�BI����b�J(f�d��"O��[�^n� �(ڍg�0e�0"O��pQ��'Oڠ�aG�9-}�27"Ofai�
�q���(u,<m�!"Op8�b-�)�&�Sa�%	?�]��"O��醁X7
і(�'�Lq:���"O`�hĩ�+
h�	$G�	N)����"O�`*tȁ�h]`�P��+�}�V"O����o>4.f�{�gB�	 ���"O��"� �8���p��Y�H��"O�|iB&ڮ+D|AAT��d5�%"OjD�4c� �N�:�#�� Y��'��	Z_�� ��Y�KxV,Z���65��B�	'	Y=Ё�O.!_��r�ʕ5�JC�	0^��@��ĢF��]���	2Z�C�I%��x
�[3):z�
4��,�C�	� �25�� A?<S��a��՘
0�C�	.��t���u����VFY2��B�;M�XYǨ�}FD�հS��B�ɗo`�E32�Wi�dT��l�9=�^B�ɽy��99�*��6�bE�4wZB䉸r���eݻB�F5iG�8>B�	 �rE� ��+i&�f(A(?B䉌.�yڳ���# �p�:�1� D�`�w@ WӲ��T�)%�t8�bl>D�܋��s��%B�H�^lx�j'D�`{�L�K�a��)J�k8deY��"D�|���&#��H����($D�X9`��)���(�̣1����ԧ&D�4aNO�\{�5�WO#q�t$Q�%D�dQ�����y�xP`��"D�0����,���c���
'�՚�E$D�`�!)]0:x� ڸH�r�Ғ�-D�x�Æycd��nU"D�pٺ�+D���I�����ԄPb�yb4�(D�L��Sd�ʽ��РvE�@(D���d� 	-�(I �A����'D��;�	���q���+Z�H�aL$D����Ø18�� s띍>h^�b	/D�D�U�d0�6I�8�������-�!�d�	L?�Q�lҭA���J1"�-l�!�	*�����������׸&�!�0��͋Ck�:/��/��`K!��W�dɘ�4,"�8��ۆ)@!��P]�P ��N0?-�E���D�Z�!�>`�BG�7x d�Is!���B��@� z~�K���[!��<f=�u꣬Ȧ&O����B�!�]�1�XTqW(A6@6�)���)"�!�� ���N9Ve2`����X�Y�"O��R��{.t�H�]�3fu9�"O^���'�;(��˦/�7<�RY �"Ohx����+x-���5�	�p�m*�"OhyЦ�ƊCعڕ��&�^q��"O�Y���2:8����鹦"O>�2�D�D  ����)���	"O���tH���� ���0� ��"Or�IF�(B4	�J� d��"O"h�@�<�Z��2Q�-w"O6�0DX�b��F��ݤX�"O,��M�3AU���eZ @�@h�5"O�e����&ˈ��V嗏���"O�[P��"Ed������9:�"O���'8^SԼAs��`�ȍR�"Ol�!�f�:��9	�b�:���"O��pΌwuN8�F �`��ayv"OZl�E �Y�B�0V�ʾ�*)"O�q��������_�X�aA"OR���ą�O�����TKT�˶"O��2f#@�I}<Q��Dӣ.�浪b"O��*��޴.�X�!���d�W"OD%�Ȑk6`�v���K�򜹗"OjE�a�3 ��ҥ��/)�≛�"O`pa`�_k�f@�i�*E[�"OnI@ "-�uxD�q�}#A"O��Y��2v(�0"�/�M��@��"OB%3C,N�~@ ��%��p��"O�i�l�U�r�ڣ,	�)�b�7"O�e���~R:Q�0��$3�[""O)�M�'j�J}�������"O��S�&�#/��9� �Xy�`�`"OTj2�W�_��ȉ1f+ZX�9&"O���A�Ƌa����vă3H¥R"O8���1J]( ����!Q����"O^0!jT�!tPs7�*( (V"O�AQG�TK��	�#��X%��"O`��q��H���$�Og� i�"Of�s+Q�@��]"tF�z�r2�D?LO��4��z�B�XSެ:���0"OP��.R	o����������#"Oȱ1�4a,]��N�1z:�B"Od���Тk�b��.�,Rh�q"O��!%g����x�t�ҵ
R�У�"O�:��ȏY��*�El'�\�"O��8Q�Y�h?�(��#\ H��8z"Or�J�^��6Dq���{�^	��
O�7-S�s�LXU͕�hU^�1�	\b!�ĝ�KUz��BJt�, 8B�sO�x��I=WVt��I�=rU�U*�T��RB䉪c�>��&�X�w�H�a��M��B�I�"[�u[�hR�D2������v��C�I�)�V���J�D���a��WnHC�I07���H!@Ҟq9!Z�{^B�I"��j�m��@4\1�@����C�I, `)��H�GV�[#��)|��C��+>�@,r���@ZZ!0��7E��C�I>J����T	�0y�Y�7.�C�I8���q`M�'�"����ۍ]��C�	�O48SFa��>�e �ك"��C�#d��D��J/��XЄ*�MNC�I�{{��c��}�\µA��K�(C䉮߾��m�9����ԣHHVC�$JuԄ�C�܆S�r��kQ�n��B�)� b4�PoT�?N�x��P�3j���c"O�l�$�6o�~ܛw�'MXd#"O���D��=�^��,Y�'��heR�<�O���$�A���s@I^�!��\��`!��3N�ℏוwR��[WBMe!�䒽�p�H��.�(а��x!��%|�������J9����0�!򤈝Y���'�'�
!A��,�!�Ĳ}��M���=��m��e��b�!��x�T�RBX-L]�X��/I��!�)#�<�P��ÃOH���/�Py�T( ר��աG-�0�J��P��'eў����ʑ�B2�2R��]�6y3�"O��ꄬE	2t9� Y~�p� "O�����=\�z��$�A.;Ҽ���"O���.�^~�����;yt�е"O���2�K�^Ь�b� �1T `8!"O\4�ᆊ��&؈�{@x|+b"OR	�b�;9��in64\��"O`P�l��]q���-U�8�4��"Ov�k��F��
E1t��劃"O�(t�M�l}	 V  ��"OČ����H���OM�X�a""O�8�D�i'��!���XU��T"O�u:gF��~��֤�g�
���"O� ���	�Z@�`�%Ձ)Ҩ��"O�\��͗!� +#ށS`v���"O�L�vGM�ݖ9`1G��Z8ؙb�"On����ի#�0��p����l|�7"O�Q'�����CƐ�벼�p"O�g�K�9�����Li�"O�M��DU��Y�sBU�=��i1�"O"d�AFM�08����ܡ��Y1E"O�����vT,Q���"P����"O�	�3��E8ڸѵ�ڜ=y�4@�"O<�S$c�Z��	�đ|\:�kw�'��D��($���y�V]�fh	�<v�|1��+D���qD�;Z��(H�w�x���6D�|��L�IXZa	t&�8�,��4D��#���z�8���� PQ��a�.D�$�T+��2�Ĭ�d� R�a`�(D��3��02ԳshT$b-�P��9D�DҦ�L�d�t�ddS�E�~�ZD�1D��1�I'hj�9@�g&���!,D����όVJ���E�	�BP���)D��A�yO �@�e�z��"*,D�L!�؋8E zq䓡+���,(D�T*�"�@ IRֆ�0�ʒh&D��*�%�6��ASЉ�8o��P�?D�tc�韂p�]���<zJ��P�%;LO��l ��17�x0��}���¯6D�x�B�ޟv�b���'��[:�t��D*��W؞ �QJ��.Kv)��]�8XH�1"O@�ᕡ��"� w��!`�4D"Oh�H��j�����`-rj�F�d;lOD��OM�mޮ�0厓=���a"O&�%��:�n����H�j@Ƚ�A"O,�S�a�-�1&�ϻ+(�]i"O�� ���Ku$�9� G�;"�X\�lD{��)Q?fzf|K`��{��%KP
�-�!�$@�&�]J�$�%+��˵M�!��L�|4<�%��9?~��W��,=�!�DY�:� u���%<h������!���+j�3��%�┊�
�
x!�� ,��@�U�$�{�B�u~�:��'|�'4��!@��#h�65��l��%o����'J��[e�Xl�Z�*K���I����!�X��OO*�6� �-�6���"O^X�P/��;$L0y���<V$J��	b����#C���#���_�ai�j	�m|"C�	�*�ڶ�n��� A��>�B�I�w���BP�ق Vi0��8�C�IM�ޠ(�������R��C�	1AV�c4H�
_X�l�V�O�YLC�	!LpT8{��V+�L�㎖&�(��0�ρ�{�v�Ad��D�9�H=�O:ʓ�?�l����A+�>>0�ɲv��O�<q�k��t	��%�>�4x2��VT�'2ax��%OV�!2˒�zwԜI�E���y"-N�A ��
	�mp�� �R��O���b�D��O���WO(h��5��+�(R". �g"OB�����:4䬑����� X �1�O���C�U�4B��P%�<����XY�qO��=%?yۆO��:)�� hX�=,�]4�0D��za��#j�<��k[87��0�,D��(1K<jX10�.T��Sw�0�xm�A�L���J(VEYרÙfD�B�	�-�&	 �KP�p�؝��"���C䉻[��I�7C��3�ŐA&[�(�C�I��t4����X-���^���ON�=�}��g�6s���k۳�
t�)EL�<rC�Txy�C�5�L�!�E�<��fT�������'PǲUS''K�<)�NܷMe�ݑ��Jo;2$�G�'oa���&�pqݸF�JM�`+�8%e!�d�&�L"�$�i�Z��$N8A�!��%�t����:����<M!�d^p8��c�B�yuz�aW�0B!���Zt, �b�ĈL^�a:墉1x:!�3'�Э@uAE&D��@�H�!�$�n�{���L7hٙ�B�0!�D�&Ń��q-"Qp�
:xz!�D	"+��1���0m��Q� Dj!���[���,��R��vS�;!�D$�V9�0'΢6�رۧ-!�d� O�:4�ħN�	�>T�U�An!�d�O��w��H�d]��ޮ`
!򄆅6�&X� �R�,��ȳql/~!�������bF(CQr�J%E�|�!�D[� �����DǩG	�-�SƇ�t�!��P�<H2�Ѫ|Fp3qI�U�!��ج��4/\�)SK�L�%(!򄔾<�N��_����e��q�!�-F���)�M�C��	BÄ
 aG!�F��T����8����N ��ȓyY��K0G�91�HU� D��ɅȓT��!�K-F�X�c� �4�@��ȓo�@ᚦ"I?ǂ�ㆇ_"cmz	�ȓ!����D�6`�l��
u)t\��4h��$μu�~S� S�$�ȓb�����=%d�"�!=`t�ȓ4X���L�嫓엄g�>������)q��?C����#�ʸ՜t��	�I���̲{S��	㡟�U�"Ɇ�h.���
�Kn�R�	�`�����2�*��w`
'2�>�@&GM�s�왆�+K� �R��k�a2�HO�X�"%��d�&�P�F�"F��b��]�U�i��S�? :������n��%�ε#t|�q�"Oĥ)$IQ!	�B`�A$(�,�r�"OD����c��M2�f��:���8�"O���	v�����	=DUv�"O��b����H�X1CE��xA��"O-��g%#)Ad��\��C"O�04DֽxpD���E[v]
"Oh-*#��`9�9��'H�!kV\A�"O��r�M�%昍�R�� \`T�I!"O����rIڗO�^�	�&�y���`�|!"�����H�Ņ:�y�$L�31\d���O�+4��8�o\/�y2&@�{��4St��>qb�(��T��y�@@P񭎢 �h84�[��y�o_�u$�al��@DD���\��!�ˑ6�@(� �� �+��\=!�d�SҤ�g��!
��K��,�!�K?X=
�,9�<y�R6sj���'��U�E�o�b���Ɣ6E��{�'
Cs"J�#��*������K�'c���ad�92+R\�S�M�\*p���'g�Y�T�f�d��f�3>��'�X+b/�h4ջ�d�&e��'i� �O	h��P �� �.�D��'���ǀ\����SE՟2�L��'��v�Q8�tdP�J�bp*���'5�iS*Ⱦ^�0yK�j�Xk��A�'*v�s��S� ��D�YP^��'���%O�u 
���텤F��()�'�>L���4��*v����'{�$:v�^�V6����9u/�x�'�^H�q����M��%6?itAs
�'4��O�H�d�I��Kg�ٺ
�'��y@�H$t����ldD���'! �;�,_�i��0��%&u�rI�	�'��Q��CF	�������c]�$��'���kg�Ϗf�-;�Y^`t���'6I��)W1?�P�Qm�3K�ƈ:�'F�뤯�,f��u�ЩE��l1�'k��b�۬;�6p�J6Z��'X��a��A��P#b�0
 ��'�l�X�MξP��-��J �8Sxx��'�}2f.�0``Le��!W�*@2� 	�'m��:��D�1���@��M>*��ܡ�'���9ʒ#nK�8j��Q�(qr��'J��PR
�D�N�JAj�y�'-~���W"Wo"	��j�yQ��
�'^!���"�pP�3��x�&�	�'�XL����:�};f��E�$�	�'��,�r�R�kdoB_K���=D��#u�%C�-�V%�m�}�C;D�d��'On>f���.�j礰1��;D��Ç%��y��`�CN�+`w��{1�;D���mKVdFPr\N���;wF;D� ��$�r9���>:�YX1!9D��9��3�F����֒=t��R9D�H�C�,b�H����'Q�L%��!D��Yb��?�>`чM�0~BI�aK?D�\��i@=��8�H�4A5
<D�ty��Z�V�M�NQ*��aQBf:D�,�f��A�.Q���+'����p+#D�db��p��q㏶P/��p".;D� A����,Р@��u�v��,D�P�S��7���X1�ڣ@����7D�� ��HB+I�u�����@�O��婇"O>�	df�)T ()�i>:���a�"OD	"��P6���HH����"O�`"����7�$ ��	M&~� "O���L�u$^��G�y�q��"O��aFZ>T�pщ���ML�Y��"O~I�S��fED��-����"O�7����Ј�k�4�`�s"O�d�Q��_\���ܘ d�y+"O�q� �G�ZuA3��iH8QS�"O�r���
b�1�Í�.(����"OI`�BR�d�f}Q�D�	��@�G"O�0#���8�b��^�*�j�7"O�L����j�$�݌�a�͏C�<��2Rl$���B5�:e��C�<9�$Ɵ@*(
f�\,Km���+~�<y�6,C�����٠t� l�$�x�<�d��0<TDU���yЭ	�au�<�GlV�d��h�n�NB�+�k�H�<���� u���w���"?�T�Ƣ�E�<P�)�̅���O98��tɋA�<Q��H�6��<qf�´PEj�ZS�^}�<1ֈ��-n"��W`R/7����${�<��H�84�<)
��	�b���e��v�<�����.,��
+Ml���j�o�<�3��d��ɫw��1-�e�ֵ<B�;cH��$D�S����GLC��c���1�\閥�`���DC��#�X	E�;9z�AF]JnC��7u�$[FH!R�O2�<C䉵^�^$SF�!0��!�:C�-A�x|�įQ�\$��VN	�C�	 |��1o�(�L� ɛ7c��B�ɤ9���u@�'F����B-6e�B�ɻ/���f/Q.{u���
�*?�B�I�$nR�h�Jf���O#(]tB䉝h։z�ER�UJ����)�QNJB䉂,�Z챦E 0�	�B%V+�B�I��؈�DIM֘�R@X�.�:B�	�w�6�1c�Q l��*�;�4B�I��B]ң�O�<>���[?=�B�*|a�mĢabj�����i��C�	�L�8�D.�"S8���Y*uͺC�I�"t��`)�K��iןV�C�8����&�x�
H1U|�C�IuF<I�q�G�?��ԻK�!�C�	
@,J书h�d���'�K�3�bC䉃{y�;��?�h��̊30v.C�	M �xtN���U�vl��a�C����A����pw�}%��
�B�	�$X����<9L
5BźPS�B�I(��
W�ԫ]i>|i�^�h��B�	XV�0f�tu�*3M#��B�ɑ?�D����Se
�{A�֨!�LC��%Db4�+#I�o�>q"a٨'>NC�PJd���_2M���Kw�T)k�C�	
'yԱ;W�=7�i(�#��s��B�	�
v���4DݷI�楂'a�,rv�B�ɹa9�`C�I�/#N&}��i��&C�I�p���"�]�6�$� S!�
}�����#��ѩ@>�#���{�dS#'%�!�d����1�:h����G�)�!��96�<����
M�d�%�).�!�Dվ(wJ1;���+8��t �Ƙ�^�!�� 
89�� %]�W�J)ko\Y�"O(��@�ؤP���a���܂b"OlPΈ�BH��� =Ѻ���"OB������,`���GW�JW Ts"O�rd� �0��� 6��,Xg�Ya"O��P�Í�5"u�������3�"O@���c�r٘vǃ�z��"O<<��ㅴP�2�y�T�n�d�"O:� $��pڄ�&�M��c�"O�ء4�Z2Eg���d�PڬBq"O��A+I�%���	$�C����"O���Ј�|ƴh�+E6j�8�"O|�;�)�6��!�q`�cɊH��"O�`�Aվ6�rl�fO��Ҩ��"OLe�N�?�|�Qb`#=�0�e"O�@q��+n��U���#W�.x��"O�:�ϴu�ј`��8���"O����	�Zf�۴$�\�['"Od�����A̔�/s�Z�"O�!�@W^�<j��= M�t"OF��@�V�i��,�)M�xո�"On�H�f*^�8ɡ헊s`AC5"O$�BȆ)#�BkK?�D(6"O ��3�B�>]�B���>I��"Onq�-��r�* �_�́7"O؝�B-�?�P �eq�B�ɓ"O�,��lM�C%����cS(z 5S"OF�j��;s�6{QI�+mȊ]��"OT��f���c�Tps��͂W��lQ�"O� �ڦo��%��U��Q"O7c�BW��`�,XЪu��"O �A���6D����4<���#�"OHcC��6v���ခ�n��&"O�x���I��.X7J�% ��Id"O���~l�����-0Z�""OH}CT�������h�Z�@�*On ��LJs�N)sc%ř]� �'���3�X2u(�@�-�>Q�Q;�'5��c�.�=8rD	:@�Q�i]�z
�'�����L���I�IéM����'�ta`�'ݶI�d��ơNrL���'���J�Ɏ�NB���Vj�h����'�L�;R��;\�\%� Q�k�����'�h bEh@�|ip��:o�:A�
�'����J2Fb��
 � g�`e��'�1���?��X3��U�eI�Iy�'|da��h\lq��Cҽd�8�y��'6Z��S�^�r��Ї�
�Y�r�x�'��lɱ�}�ְ����@�&��'��-ZU ���2��Ց���d�<�&�=w~͋e$�6�顱#�T�<�&�[>R̠
��JX�u��@�h�<Y7��~��jVo_m��`�E*d�<���2m.6���l�	7l]aF+^�<��9�\;���3�b��%�D�T���C�(��iڥP�,m�����&��ȓY�` �%��4���9�Ǔ�5
���ȓg�аr��!�8��R�Y�Fen��ȓ7���:⥉�q���H��T!M@0p�ȓ,I�m�"��+K|����]�$��ȓ"��	��C0$��hBn��Q�t���1
b��#��M��ufK�o�px��]T�a ��r��"
̶Vʂ4�ȓx}���bM*�� ��� ��p��S�? T9V�j: ��r�>Jɔ�+�"O�=Ө31h���>	M�A0`"O6���$X&;Ӝ��a�RB�Ikg"Ozd8�I�9��x�m�;6* "�"Of�In`��R�m�tGj`y#"Of�a��XtV�	:.O�\��x��"Ol5�Q/� n��� �u�4���"O����{�����I�d c"Ofmɗ��
d蜫�"_28ھ1�2"O�q L��DP#�� V+<�2�"OܹP�����q��A�a&�,�e"O.�['�&���K�H��!��p7"O~A!��V�8$�@J�Ƽ��"O$��T%x0�	��+V�"y`�"O <�7�P�jo�Q����t�T��a"O�"ɲBoH+"G�8a�j��"OT��&�%<a�hYƀ0�d�"Oj��w����Yo��{�HA �D0|O�hElH*A�y��Nܫ1�=R�"O���ÔZ���kA)&�4��"ORL��!Lc�X�F�<!�$V"O���ϫ`h�%�A74�=��"OL��)�?"�d}�n�=	,d�e"O,��Te��b�V�(�ҍi�tJ3"O�A¦������ǱD�4�I�����E�$hݜtP�ӤND�Op
,脣��y�6)* l�'�²7���k���y�o]-	V�ٴ��/���	��y�N�'�D82���(iQb$;�y� u���`A�֨$w�Y� o���y���D/e���/#�H{0-S�yBJ�$_P���@�71@��W�_���O�˓��O�lx��S+IH�M��4}L��I�'t��bQR���Af*q�'������X�td ��`�53֜[	�';�"T�j��P�%��2B�'C�-��	�n���S�&��ԋ�'���)'"����P�/1�����'���]�F�h�QÃ@'4ݛ����O��D0��u�r	㖨��p��F�\��B�I=LS$���m��ؔp	��w�B�I#g���3#�0<�r�k��	(r �C�I'\�P�NNu ���Fë	�vC��F��E�u�0��Ъ�m��"B�	vVځB�R(�����9m�C��*;���;�$�Nd��"�.;�C�	)B�$���D����7	� \+""O>ě����j�SFG#��y
�"O�h�G��U��E�Y�d�:Acr"O*(qԄ�����瀑��q�"O�Q5��$-'>0jS�@�z��qpR"O(���B�:�0�L��t��t�s�'�'C�%#��>j�`$Z�Iۃ<e����'�ў"~���Wr�T�ȱ-D�9���J�<�B�?(F��&Ӣ<�T����C�<��MJ����e�|Wތ�,Ut�<QV�׳0vbr�)$\�A�As�<A�IT
P��ȊU�K�9<rx��bYo�<!#T>:#����B��{�|�؃F]V�<q3����4�I-D�403DH�<��D2$�R����>s�r���(CD�<� @l����8�d��a�}�<qwf��(l!t�	�a�>���m�C�<��ɢ:��e9�Ț�C��B��h�<� �ha���8fj��8t����;�"OX��l�
{܆L�J�0���[C"Oʕ �Oɤ;������G��ؤ�A��`�O�P��֧��5n��cR�H0�`�B�'gp���ۛ+�}����'����'���Z��:RX|�bˑ=0k	��'���R^*�Y�)՜^���A�'P�Hq'��]����c�4^F��	�'���օ�7�jP�Q�I]�F��'�^)�)@�-�zYCD+5||9��,�S��KۮT��9�(?<rZ���Cə�y"�G �h� �&�,>ڊ�z��yB�\:�beL1Ehj��EMK��ybOU�@J嘐���P��X��M1�yBC�4�.pr����Fr���E
�y��V�V3��:��Y�Bh%;��4�yB�Τ/\J9�F�Г:lQ"VD2�y򄞍C���V���5)R�ru����y�Ǘ20��R���yD8�@��y2��#Dz��X�9v8Yaힶ�yr^ K] �H�M�68JFd#�I�y, !TC�`xc L�#��PSW"J0�y⫍�HU���ꙴ!"p�Xq�_��y�D�*rTɣ��޲�	;�.AIyў"~Γ_����ݭ2v( ؑg=	�<��	���5�R�3��U�A6 E�ͅ�0tl�9���p@>9�E��/CJ�لȓl�nٺ��D�Gu�P��o�*��P��D�M*VF˂d�mYu��+�$��ȓu�&]�Qe�{�����y`t݄ȓy��I"�$N����E!�f��h��SVT�	� �Mʚ�$�dd��M<�����s8t���M��D��0&����*^����b 	� 8������w	0(�1A�U� ����E�"$M�{�J9 �利��Y�ȓu]b��!�PE�� �^1��؇ȓ:���C1�����f:����v���˚�-f���G!\>oU����ss�8�%M�z	����+�F6U�ȓ�)��C�-
F�����&sxd-��8�T��Pn�WIJ����y��Ѕȓs��`�'e� ��t������,����j4*=��S�԰r���ȓ
ۚ��t�.}D�rꀪZ� p�ȓhv��q�Ú�%���O�PW�U��pk"��a�E�D���1���,%>���$�h��+�� 8v�9é^8;����0�ى6)+)6��V �;\T��r(���hG�m4�h��G�+J��ȓu9B�a�J1A5�-2!шX�T��ȓ�౒Q(�:���aA�Z�mB���P��l��� ��g�豠�,ؘ���"P �ȓJD>>�0q�\��腄ȓY7�L��"=�0�����{�*u��2j���Q7�f����� y"1�ȓK�u�!�q��iC�&�� �$���6ƈ�8v�����w�P0* n��ȓ+���͟�Y
g*ݐު �ȓv�4�ˎ�#�~�����O l��JD�����4P�\�����?��Ņ��*5ːIS���qy%m���ȓR���Dƅ�Mf��.�1O�|�ȓ�v<X�ǃ�w�(M�`f��:�f���S�? ��S�D4>��u%Jr4�c$"O	�,t D`�I�x�� �!6O�D!�)�'n�c�D{�p� �攦j�bm���:yH�EX�>>Lʆi��F�$��tC��p�lFx��0@'&�Մȓ�*��*�	�� y'�ݞ(-2i����A��G^�Pp �5e�H\�ȓ=Y���vW>��e��3*�Fl��"O`(�af�uan!r���X�"O�9sb��xg�yB��r�h9"�"ONL��Lր�`�s�Ј�N1"O��)�%J	h�8c��� ͌�H�*O�ఠi�	�v����9Yv����'H0��gߡU> 0-U$�ܹ�'����Fi����` ��
�v)�'�;��
wIN�c!	Q�qEf�	���W�����L(T��� =����@���"��,.(��+b��3l1�m�ȓ	����#M�_��CGJ�1V��,���r�ڞ :� ʕ��t�x@�ȓ-?Y�ट<!�AB��[�d��f��00b�?.�H����-�`���|ڲ�°I��A+A�#�+04e�ȓR��
Gl�>.4	ѧNX�H�~���##l���f�Ҡ�a�@@:��ȓLp����L-A�zY��H����ȓ$�*q�O6w���!T��-�(��ȓF3FYp��j�r�
����І��?��$�Y���P��m*
p�p�]�<a-I;Y�$��M�O[�D��]�<9"��o$�D��~���m�\�<��蓿.E��C_'R6� ��Z�<�鋙x��W� ]2(aÏPP�<��Ǆ�P5��Z!̘[�vI �D�V�<Y�A�>��)*s4�A�u�U�<�u�_�~�ژ�g Tۄ ��T�<���=�j���V��3�E�';ў�'},�H�6�л7�90��3���ȓi�ȡ��ˠA~�0�j���$���&��AE"�(�"$&��P��M(�4���hf@��A@1��ȓ3�"xi��Mզ��$�
m6�ȓDI���0'��o��p��7Hht�ȓg��q���zK`a��,ڐ<�����"�(I�#K-U*^����L<@����nŐ=�4KD�I�ۃ���\�6h��R�l�����^�A�wF��}�����-db�[��ӄ{n`�zAn���e��4
���,N&M뵨�+�ԅ��L��3)������p�ֿs�d���
0��J�7�����,�/�e�ȓAV.�U���EQ4h�6OI4v:�D�ȓGBJ�X�@\�m~Ft� �̔!���~U�sb����XC�ީ+�x��ȓa�*��=˔��ER�b��ȓK� q�Q(JF�B0��}�Q�ȓ'랑kËƅU�d.p�ٕJ�z�<Ib�@�R��p�̥5B@9�EAt�<�UQ6G�⍢�̈""����2+�D�<Af�̴1HU�Y>��ve�<��P�L�l�G�S������w�<�S�Z�;܅�ҥ�Hkh6��u�<�w�	��YE��=+g���`�s�<9��Γ;a&�A&�84_$M[L�h�<� :���+4ȑ��,G�,h\�Kc"O=���˹f�vQA��M�^ �c�"O�X&�<E`|0憈�H�jTP%"O*d��
�S��dK��Am8튐"O���V�ޓB�f�yB�O�z~��"O�!i�]�P]j��E4:ef��"O�u���DaLP����&:/~���"O�]ѱ��(<N܍)T�OV���;g"O����JR�-4tM"ԉ�D����T"O���^?/�d�yF)�1 �D�d"O����F�-$P�N��@��R6"O�8c����B�H٦,�!���7"O��9w�^�FK44����3"O�xB��->��0��)���"O@�q0ǀ��*���J%"����"ObT�&̆��M#�KɩF��}1�"O�thT��0Q���2�K:,%	�"O���&�]�	��|swj��n( "O�t��(� ���d�<�\aZ�"O��`ꐔ(W�=�Fl�."�l�� "O|X��H�;��ls!��/��hQ"O`(30�"�{DjM�k�z��"OԨ{�n�;�j�Bj�.3��@��"O���'A�5����: Vl#"O�d�X? ��d��&��i��"O�h��޵zt^Q�T$��G�M��"O���q�!=��:q�ƀDDQ9�"O��e�%��p2��*\�nme"O�QҁCD����7�X�""O�A���45����F+2�a��"O��q�FU�!C� Iw�$n1�8s0"O�$���ʋu���i���i�f��G"O�q�UHݓ:ef`���T� "O��c�I4�9�tF�R�j�"O��g�X#�Z�QSo�48e�Q"O���b�ۆ>��cf�B?�B��V"O�AfJ��^Ȉ���^o�Dh�"O�9P�����b��ոG"O�E�ՂM#������޸H,��P"O�L[sjݴ_<Ph���3%3#"O.Ջ�X$D*��y��V�Z9ۗ"OZ��� ��B�p��^]O��A�"O$�S�mɰi��;��1�L5��"O�"��ߴ2*��6�JP�t�Z�"O�$�m�'�|�2cF���v��4"O��[� �$=�@��X���	d"O<@P@�� ,>$x��y�\!"O�2��[�o"	�Pd�]z���"O�Q5� :yvx���	�B_0e�B"O�=y2b� &ۮ�8�ʬgl$Qc"O�t!`D̊0�t�Br�2
|��S1"Of��2g�
 ̻�*�Ot��IC"O�UC��Ų}��w˝ci�h�"O��b�0 �����At4!��"O� s���f�բ�ԧ!��	"O�5�N��88WJ��fo�t�1"O��9�J
�0dS�O :
��5�6��؟"|�'Bd��"Ǔ)	�I��*4�a�
�'�ri���7?.p�S��)�P]c
�'s�(PJ�?	L�ڵ`��$�����'�
�i�X�@C�E�bU�Q�>$��'�vi��lY�g���Z"i�H�n5Q�'	��jظ4y�"�m��ű�'v�1�SA� �q0�B�-V�­+�'~�'��)�3?� r�I�*��[ < �JW��j��"O����`QЄd(�NB�|�J�K�"Ofua��',��u���;��e�"O�Y�A�J�Z���[�8r�%"O:e�v��-��SP�]%j��1"Ov%���
��E��NM0i��pq@"Ob9���ܜF��Q;rM�&�����;�S��yҬȏys���̝_G��j�S�y�(� #�0��/��[���U�F��y��*vƩ���C.��1�d���y��סN�^9�A"�,��r#Ǉ��y���35�ؙb����{�6�`���y�bC 8t����y���
�����y��U?o� ӳ�X� 6 l�wN�y�&
�_i�Qpw+17�4���y"��1�.�h�~�x�'�-�y���$ȼy��*@{�h�)�皼�y�eՖ���9a�řzd�zկ���y�h��jT�\�Ѝ[&n�"���ֿ�yR�J=,v��#�o	�2�J�"A�8�yB*͑7 �$X� �s(��y����%d���C�$�P���yRD^<�e��E�q�p�c��ʘ�y�I#u�=�p��f/V`I�]'�y���*D�U�����o�2��y2c<Pżps�c�<0�⯆2�y�H_�;&���δh�Щ��A<�y�`�3{<���.{W�5P��O(�y��K�I� ���z�&�� ����yB�޵l2(1�m��w.���S�� �y�II�7�ܐ��n3r��LY��y�I]:(�e���_b�* �y�c��� P�X�*���tc;�y�[z���^7"f��C�͐�y���T��aa�|��[��y��1N��z���s�^}�B�y���]�)�� �3���+A�	?�y2 K�r�j$�@:~���P Ѡ�yb���g�,њ֤߆gn�$�P$'��$�S�OOh�4h_�e3|]V�jZ��	�'�h��F�;� �el�).r=�	�'~yM��Q�m��,��<��I�
�'�L�����􅰕�@ 8���	�'Lh-:Ph_�#
15��!_��'>r�)���, �Ĭ�%HX'ex����'�^�a��D���N�|��A
���S~��)�'(�p�ދ]
��$ᄉ|������	����4��Ē�Kh�ԅȓixè[ 0�4���MCf��1���j���@���R�4�:��r"Ob��1��%[�����A�'\���A"O@��ULҦ^��"���N���� "OĨ��ݱr4�I���ۙ~���3�d6�S�'Jo^�#�O5k�Hr��R�����ȓ:�H�7n�X���q򡊟c��p��!��@��Z�U�f�Q ��UwD4��D
V�8	J��&mV~x}��~t���'+F�Α
��ՇV� x��e��YC&��:���oI#Gf��ȓ#h�����Y%m�f��'�!� �ȓT��ZH��F a(�˙�g]��YGn�`��*8�����jT�i�Ԑ��*}G�g�H��q	� ^j)��Iu2%���SIR�m�P�М �����S�? l"T㊃~QF���(�y����"O�P�5+X�U�|��e��2����0"O�*�����������9�2Pa"O| �R��|�p��H?,Lƽ�"O��@1(x��¨�C@N%��"O� ¡��45��pD.H 94�q"O�!��B_@70m�A.�#vL�Ȓ"O�� �hħ;�,��ܪ9h��C"O�b��ߥt���!$���2bJ�Q"O���v�޾+�~H����X	##"O�`����8i"B(fM<�R$"O�� �	�Dʁ���'Z�
"OԬX!U�Dx��*s��b�"O���o��D�bᩙ0���"O� ����k�0�C���H�P!"Oy��MΡ=���#�"�5r|�ő�"O��1&�wD��5��ci����"O��(v⍃mRh��"\\�Lz�"OȌ9Sc
�4�
E�U.̿W�d�
P�'�'����U�a�ʄ@�^O�x���'�n9�.�5�Jy���$rR�9�'�̡b����L$�!kQoX�  ����'*����2���̋>`l5��'����S��'<@S�G�>DB���'�<���L�J�6�b�~i��'ݒ8���ځ�@�v���V/���'��<�q"QnN��e錙�����'��sL &H�0	�K��>1:�'	��MA�N��\�ê�!m��	�'Sn���ͤJ������j�s	�'�`x�1�Ք��M" ƅ> ���p�'�P9ѭ�!Eh-a�C�0E�\��'��A��S�ʼ	 h�?��k�'�ڬ���:h+� �2�[5�ԕp
�'Lb�+�f!\<&la��G� {he
�'�����DE�jɫ���!e� �
�'�P� (��RL��0�ĝM��{�'���Γ�AV�����J�ιR�'� �0K�(�f���=�8z�'^%���ֵ��C5�؁$��X�'E�	�W�6CTd+eV��Ȱ�'!hHh�F҃@r� cD�@�h��'�Z�p�H�:88ܘCh)@`�qZ�''��q��T�Q��cM�0����'vxu㭑0w��� �N@9�XS	�'���7�Z�H����E�(	���'���d�%{�T��aa:1W2���'�Z���AÎB�� �0�~O�ܺ�'}�������됄�A�j���'�����I��D�B�L���'��XAtڸ�X���nC���8��'��iqa�:0�YK�-���Q�� ��}A���+���E���4����ȓ=%t����T�P�J$0�i�#>�Х�ȓ6֜I�#ˍ�tf��{��K/b-��M^��3&J�V�*q�c�2m@)��{ϲ��M�06X,��a�>�����a���8�%^k���ę�nqU��g2xIA6Mį/x��ċǸ�!����5�eƨA&�T�Ī��Xt�����{G�Ʉ}P8@	��gQ�Ɇȓ:ў0!�&�$g��Y��C�A��l��!ͪA ��E�~y)0 ՜�t@�ȓ �0�7͎�W��9Я�/%�]��S�? ��c��
?>*�����	w���*�"Ojɚr��9A�U���	~��LC�"O�Ȳ�c�BwH
� K�Vm��:�"O�RW��\:M�f��(&N�XP�"O@����[��Zs�..M�AI�"O����*Цq�R��veI$[;�!��"O�p��W�0V�`���B��p{@"OV  3"8G�$h 2d¹���kB"ONk@&C�Q���ǃɽE<����"Ol�ʂ�߽���h���"�!x�"O�E��u���7��l���=D�t��0l�x��'/C�q��*<D������E���#��D�~K,��69D�D����E��8�ì>;��7D��A�N��a�~�k��AGTꭙ7�*D�|Ä�U4n�8���58ɨ��	#D�j�
Ip���� �Հ|���kP�-D�����Oq��@��&f�2L1�i+�OB���O�Q@�O��]����ˋc�lkQ�64�4hQ��4n� �pk�9�T�jV�2D�t1���2J�P�И�D�	t�1D��r�e�' �,`�DΟ1��R�!D�X�#�Ş)��X�'EJ3[�ݹ�5D��H 
G�*�#����A��J
2D��ɡL���Q"�D�<(����+#�O�˓	q���Ft{θ�g��5a�p1(�'_b�x�Ŗ�=^�+Sn��Y�,@�'� ]���P^X��	v�(��'�.5{�b��p�5%f�	J���'��z�%��I3��oT-����'n�<���ڶR��\�C�M�	�Y��'����VA.l�~�#��X2pp�'��	)�Jŋ��;#Ԇ(f�L���ݸF�`5Q2j�#E'��v�Ȯl0!�Fg�x+���	l�
��CD��(7!�D�()�d���9���A�h:!�K�^,����&IΆ"�)ܿF{!�d]"R8PA�/L�Z �&��{!���<���y4�Y�/>��cG�S,|�!�ɧ�}22T�>,ꬉQ�Թ�!�$C@D<�+�R& &���'��C!�$9{4�Y{5@F�"�eR
�$b!��B�FT�Hk��vM�&x3���
�'M@�p o���<��`!V�h�5��'�Ҙ��BJ�E�Н�P�U7tw���'Xh\т�x�x����sxJ3�'��y�0
Ʀ(������kc�5�S��y�I�`	\y� �פP���ybነ�X�cW��r���Y���3�yb��|eQa���k����?�y"]�4Ⲕ���k)4����y�=�5��!ҙR}��ق-��y�l��.U(F��Z=�m�7�֙�y�$K1rF-���!;��	�!C7ў"~�jel�+�s%�*P���,ג+�"O`]�$���{B4��(G�Q�hl*�"O�iQN;gX0<���T'C�0q�"O�ِU�ً��Q!�(Y+"�^ �@"O	��Gui���(4)�-ʢ�8�y�@�^h8���J"Z�n��Q����yR
F�-gaؑ�ړ#��간Z;�yC0m����l�=1ɪ1��#-�y�΍�ע�rG��J�����y*@)'�23d`J�m��k�	]�y
� �۷��u-�,�zȨQ"O­(�g�<l��b�	[�h�B "O�YÙ�ܠ���9\�H��'"O�|�F��#/��Y ��r�`X;�"O"!k��Z8X�\ �nI�B�4 �"O�pA�����q�-�u�v�	�"O&�p�)ۡ]�2\C$-�7	�dHG"O��X��@�a��Ւ��18�D��"O�Ӱ	iH�a�Y�Ls�"O��耮}4��$�2B��5�"O�ԑ�A� �[dB�޸a�D"Of�'�?g�0M���_�LI	�"O��hAl�$?���D�����"O@D��F��~K�aR!��m�v%"�"O|`�.M,�,Et���`�f�Rv"O�8h7�S�Vz(%�*_�����"O2��N+0�z���Q�X��8�"O��zu�U�+�
\���W�F���"O�|z����M�@A �f�+�Ҕ
�"O���O�#S�!{re��j���B�"OPT�&��o,���D%SE��E��"O��R�KW9c����#b����B"O�D��|~��փ����� "O��rC��9���*S-Ǽ<�l��`"O���㥞6H4|}т�����$a�"O�M)��/����J�c5�1b�"O20�f��*���)@h*B���"O�ܫ�dC�jv���gA2	D)!1"Od���	8M��9+���a3 ��"O��(�ڟ
���&��:�"O�p��m��k�z���P ���A"O���1)D�3/~�2`(G!4ld��"O������8휩��֓1�zHҁ"O���'��u�|a�*կ����"Oh�#O� ������V?Z�P��"O4��3�ХXp�q	�0Or��!"O�%����w��5Ac�\u�z���"O�`�@�@�b�,iB�&���0��"O��Q1��#:��i8q��=�*�1�"O��┮;vF8Q Gϙ=�|i�6"O��������j�&*\}r��"OZeqA^M�2���E�&t�!�"Oh%+hԍb-r� �N*<}2YB"O�)е��ƅ�3�Ā>�N`��"Oh-K�ԺD�5�g ͗".*}qv"O^��qC�%yjЍ�W�;��ˡ"O6��B��	��X��$U�,�5c@"O�	�@k��p���#M Z�c"O~����6�ě ��2I�P�"Ot`��'Z�JEqdƞ(�z�"O>���11jb�f�!��E`�"O����ĥIB����S�$-K�"O�	S�ō�n��JDg���Jg"O�0�TM�:y��9�������#�"O��0�0Wh�*!� #�%�F"OB)H�#�c����C��=�6�`"O@��cg�n,9(�A')2��R"O�m+q�2v�P���R1M�|�z�"O(sc�+_�\x�Eї(�z�x"O<
@�~P��z�5��rb"O���@ą��#I��L���HQ!�D�Q4�d%#Z�>��W[�IF!�d�;*�^�(7��W�}r�0V!�w�"6�v㤜;�E^"?!�� �h˒iЂ-�<`:�-B�_;X��t"O�T"��'��8�K];��B�"OV�Q'��" �P�j�-
VL��"O�hrӧZ�D�)`"`іH��yJ4"O�=KQ���`&l�1���Y��%�#"O�|��#n/������9M	�"O�\J*._~�� �N��)�"O�1���DH�fU �����"O�5ZE����N�#%��`��y"O�xKe!نU i�N˄o�z)*`"O��ӡ�ЩD ��*�$�zb"O" ���̉o+��'q�d=[�"O4���P��1��BԞM���W"O�8���٫*UIa�̽i���"Ox��IĈ>D�ҥ�I@��`2G"Oh{$�ύIT�S�G�k���Z5"OƨI��ir�|ɂF�����B"Op��tJø@�TcC%�<3��k"O��@���zaȠD��/,�P&"O�J�G�]c�1��A�8a�p&"O��[q��$w� �TB��E=�u"O6��e_!A8����#�1;�]
�"O.�� �':'����aR�~�.��"O>�[Ė"L ,
��,N�F}J!"OL��=<�L���*�R��"O*��cW�6Nh�c2�݀�H5h�"O��A�,4A�h�I�C9	2 31"ON�$�\ߚ7-L� �����8D��ф�ҿz9Hd#��;or4P�0J;D�\��/ϩB�P�à���m�8A0M4D��0��$,$\��Ɵ?&���k2D�;��J[�\��&���$�a/D��S"؇��y8nڀP�𫳁'D� �pm ~��uB��%X�ެPf'D��fc��%�HA��2*b�P�T�&D��3Q&�}.52�A�.	�Dk��0D�$I&��_���y��G�D���Ѕ.D���R�[�QwJm�`" �B��õ�,D���˳I�L�Ze�щP��ᰁ	5D��cR�˹B`��@C�56}L1b�'D����hI�ff�a�JL9I>�9�+'D�|B e4K��y�&�(f>`�0��&D�H��`ؑ��P�m
�}6&B�2D��␢?|3��VlI�X�ZM�a=D����@�K�|X��iH�D]\�rĥ;D�@AA��d�XZ�-Z*�t��,D�����k���hQəb�h���!+D���$Ȟ����I� �"�D�W�)D���lɮY�"��~�4 �a`&D���tJ,
�8����_ht�t�$D����Bۧ]Ė�!�\(0�$J�J/D�qp���
�1e�[�@���S1/8D��8��(��USE�-D5�q�rc4D�@��*��Խz�U;lNN=��5D�(��@�+���{�/�0x�Z7�.D��I��Jqpz����3ˌ4��*D�q��� q-8�ye
�2lqd.;D�<�F��
XT�0��� b�n) �7D���$��HPD�:t@�YEN2D��I�j�l�z��$��58�v�h$D�h1q��~x�(f��N�>uuD%D�Da%Mܞ8�jS0��g���U/(D��{� �=2��Ñė-B��Xbv�*D��lE�Wu�}9�dP�>��L�L;D�� V$9��;{���7�Ρb����E"O����ĕ'&��!���`���6"O�4;�f��[B"�Qk�4��h�"O��DމiD�]����"p"O 8�0Ȍ�i
��W�F�?����"O� Yo��YZ �ڀr4�I��"O���gH� Ѧ�!fT�$,8zd"O�q!����c��3VSdf6�0�"O(<�S�B�*XZ���rI$�3�"O�d��FA��a�G�F0t���`&D������/�&	;��^h,+��>D��9C��&��[�/�	�x|ѓA D��PL�Q���T-�P'@D"�k>D��(��,o�\жH�57�"��<D��Q�cG5;�T<�V-�H$��=D�cG� (��HՋ�;'��	[�8D�\`#�B�Y�g[u���ʦ�6D��jr�MT�:���׵>�zx?D�T#�-���<:f�-ZLb�J;D�ȉ� ��P�4�T;E���*cL$D�<(�H?D
|�2 쓘$�N���($D�<{��-�<r���4]hD��&0D�tx���k��Qq�(�*�B����0D�P���dmz���aEj���"D�l�w�>gf(�1��h�bq�3D��+ .��BTi�p���;�1D�XK���8:�����`�|��6#1D�p���J�v9>�+��įHv�lyTl2D�,�5/��t_�p(wF�\��1D��i���0$�|]Hw���}��ؠ��3D��P�M�H9��K�}L���.D�X:�`�}�L�ύ��%J�%+D��5ܪx�p�eÍ�	}�kV�*D��9�˗�yR���,�;w��Sgk-D���R����d�s�@�%Sȭ�G�8D�92�%��I�'�Q�	�V��6D�|���>y� ��� ��|yE	7D�XZ��Y�>{�l�T��'�%ѷ�6D�$˒��+[�P�ЫR�ؔ�y6�!D� �&B�|O�<��^������:D��Zp앉8s�M�����gʜ(���8D�� �h��Ib��swO�&u���%!�D7���B��J�5��`q���h!�*�^�r+��8���Gk�1_!���4v�)���`��T�T1,!�dC9(v)b���1��!E ��!�6?����K��H��uc�!td!򤀸R��Y�ͅ1�X���AH�_]!�Ğ��5rpƀ y�p�`s�>!��l���Ŏ##v��D��;�	y	�'�6dCU���I���ɤ�!��T��'fvd+O�(dO��v�@
B!��'Z�}��_�ZO��(�w`�Б�'�<�k���K�x1e�� m�>0��'��Q"�$_��lڔ�J�c�<"
�''aH��ބ V������3쬈�ʓC� �Y�y|mCe��"RD�ȓr�Nt�󨂴	�z��e�;6�P(��[Z����ńx��䠢G�6�.YDx��'bHS�l�(i��,3c�\�8��ߓ�'gd����+ }� ��X�����'ji��+ɸzŚ�CU}H���'T<�Q��ȶ=Oi���#I�0�ȓ�`3C��3#�v��3mۛ<r�ː�)��� �Y[��	m>�	åM*-^�� 7"O��"��$�T���A�B;r`zu�xB�'�@a�p����"5e@7�쉈�'U�%H�Ȋ,�ʡ��H��W	���'�:5�턳hO���V.N�P;��hOv�$҇T�Բ�+D4�c1"O����ӽT�-�� ӕk�)��>a���)�!,�H�@	|��8��aO<E!��M Y9x�S�Iz�,��r`_�Y8�'�a|� W�4�rI�t�4`�7A��?��'� =� L��䄪�#ǯ\>\e��'��L�W!J�
�!��Z�~Î��.�'=�|6�*/`�lA�R��	�'K�����P���<v� ��'�B�C#�E6L��Q���"\�L0�'V��Sh�*����CO.Lxl��:,O\��s �E���Ygݡl��}S�"O��"�o]T�����-
 �"O��s�B��\zB�M�-P�h�"OX���)�+`�����G�\4��5"O�(�@,��Z�N��e�,�p"O����dHQ����@k��P���b"O�ʷL��lwBI�@���\�`	@R�t�t�'��ǔ�?)�\��ROT=	�'�T�poķ)?�u�N�y�$X�'��<���_#}�q��cS q��Tӊ�:�S��'�6���9�*H6�>��q�:�y2��~�0U ��H,)*"� Q�^��y� ��:vj��5�R+�ĕ�妒��y����"9�朲B���٣���y���"H&)�l�$>�b���JH��y��	a�z��1�H�:B ���.N��y��Ӈ%�8D; %V�/2�9I����y�ρ#o�.�HT [�'I.�Ҵ��y�n�A���:�C��X��7���yb�1�B<�I��u@�F	�y2
 ~qB���jN�<=ذR�d���'Y�{r�i7�	'R!7c0�$$�x�'X�e3�e��\1��X�Ĝ�C�P�2�'ev��(�Mf���-ܗ6�:���䟠z�>= C$M<-dݠ�L��n��W!'D�(i�SQdd����O�4��`#D�����;t�Z�W��`sЩ!D�l`�f�:�x녁�S�T�� j:D�����go�k��B
&��T��-D��T*~U�A�����o��Aѳ�,D��`�l�;W|��!#§;X��)+D�,��G@�(�y�gA�@pU� ,D�XK��T�Be��:ҩJ�mE�d�f�(D�3�Y���
�R�GУ�2D��G� �*�P摽 ��%/��,�O���d��0�Pl�5V�A�����'L��I/:F$�a@�|u�h�R�$7!��!�d�x���&��@�75!��K�q�љūǆI��)���J�E�d)�O�A�!6~9��ʢ��:9IfT�w"O�;0�L�Q��'U)4^��!"O�<���5 �,��p!��@�,`�4"O0c�"]u*�ʆM%�\`��"O����bG3 ������7��	
�'�b���E	�,�PW'�UX	�'�P7�޴9�x��v((5�04��'7�As��F7J��ӧ�z���{���'2 `g��K�,B���y��\ ��� ,1���&�,#�<�:)XQ"OZ@�� @8��0����9$��"O~dE@
?��D15*���H4ҥ"O� c��%Caʔ���@.h�|D���	z�OkR�z̉�F|I	teN+;�V��'zR�R�M��Xd|ؒ���.�(��-O&ɋ�$(ʧ%����F/���8c$��R=�ȓE�Rh�%��r�(�u5�'�܇�I�Q�r�Zv�]�~m gD)�^C�	/�v,���̹l�^��e�L2C�	�ʜԐ� ��C�4%
�J�2p��B䉆M�ҨhS��O�,�b���9th�B�[��I���K�}�x�M�1TR�?����О~�Z�R�D�.T����e,�!���d�������*{=�=��h!���.l� ��O��P
��@!�D�`
��b`�4G;J���BMQ!����u��e�Z,|	���U�Q��E{*��S��^�D� %�7A����h"OF� �~��yx �$R�.�����>�S��0Z��x�K�/I���zW#�r�~��$�c~"�ʹ���q�E1,>�P\��ȓ��,�! ��rYP˝)I��FyR�*�� t��i�7�v���"���b"Ov����++$N�Ca�B���8T�i�ў���O���Q�^X�IBl���:X�"Ot͘� �8��!���s�b��FE�����$iJ��I�B�aZU���y��%LX���
�Q
Ra�s�+�y��'��h���R�F�H�e��gdp�㓼� 
.)bϥ �Ԁ��i-r�x}%���ɢ<�����٤s��<��@)��T͓��B��5�����8`r!ѕ.ɪa�Yx����yr&_g����qȂ� �<�"��&���Ħ���,��-�S�<q�Ĝ; ���f��w�L���Q��yL�Sz�y����q����P����3u�x��i���?�'�����HP0J��D����Gh!s	�'��LI�l	�R�I��YC6�J�N'D������ *���'V[��piR%��D���'eM�=�g���"3�5����i@(���uz
QK��]*�� O�#�eFx"�'۾D���N�=ˀJƺ$��3�'��8c����(JRY�/��
�L��'���9��ڸ#T���'�4q�u	�'?p��0",�!�`N��ih
�'�Y�@k��z�ؑ)P��/?�1�	�'j�YW���V�
@���؋z�|�{	�'��}��A
�o�sө�.f�@�*	�'K4����ϭ!�nĘ���1�$��',A�4���!�5�Ga�WH����'vh��_�-�vɣ��C�TW��'�l#DOѓ\!��2穘�M����'Kl�U:S��PQ7(��|X�'Rt�!���B*��a��g���'u��aQm��,�.�� �آb�.:	�'Xv����gQ1�l�>-��| 	�'|�9Ȁ��9'�
�H�	Z�� 	�'����K@�:�̌�� =5ꕐ�'��O�A���*�f���}�C䉵>xdA��`]/JX�G
�4l��C�I�c��H����8"�8��S/sX�C�	����&ΪdZ�
6-��C䉣(�Td�bl�|ڴ��9�B�ɮE%�8;%)�^��;G�Z�:9�B�)� *���ΗF��[�`�#�d0r�"O��`>t��zEM�3�f��`"Or-"�)��� !-��&�"O��@���V�\�+-1	�ty�'"OX�h)UFxq��@�o�BA��"O�<r�K��;���j2,�i�(��C"O0(�d�RcT��I*z�92�"O�3�d�G��]+�(�?��̙�"O�	��ӯ
�LZhʤ�"OȈ�FÆB,�0�$y&"OL-m�%.׎1�cė	8��Q�"O,y#S*+���مc853��p3"O6tr��\���ZBZ<}ʎ=c"O�\:��MG�`�aIA�v���"O&Q��� �@�T#c�\�=���E"O:�����'�9�Q�Qx��"O&,�҈�/N���R��-l�\�"O��IU��y�4	�胜S���"ON��!�19M�`��%3��ؑp"O��dS,W���҆�{�@`"O�Y3Jب9�(`pe�}���"OJ26f�'I�h��a�l
��"O��G���,F:���e&���9�"O�#�(��8U���ʈD̦	"O�T9wB��e�4<�Pʛ Ȱ��5"O��z�(��3�@<�nO��\ؐ�"O�%z	�*`K��@�f�#�4Ȉ2"O`���a<N���g�<@#"O*��Ge�:���fԜ�p��V"O��1��V	PX�� �dT����C�"O@	qK��2j������r� ��"O�X��G.@&*�����!u�-��"Ov-�`�K�&�Nt ���o��b"O��ՎQ0v�>e�v��dZ�왴"O*1y�*�Q6"D;�"�:0��xp"O�]�"�̓3��\�0g��ss�}S�"O�mA�e׭xuh�����;X=�f"ODX�#��-��xq���� "Oz��AIQ)U��1���`�Th��"O�%�U�;YИ�4A�6mҲ"O)Aq��=[�@�-7Pݘ4"O�a��!k��8Co���A�"O���p�'��lh�䚞&�
���"O>$�Ԏ�� ��m;�dD�A�h\+d"O�HP��3T�<#U.!4�T�`"O(%���\a?�P�6k�6^�<9c"O�$1�AR�,դ�v��7f��:D"O(�:D�

��A�)D�?��`�"O�D;�3f��ЈY}�P	�""O�l�"�ӭ*Ԍ�js���l��!���'��'8g�DH��@)��!C�lC1�!��,pJd��/=���؅�̦,�!�䄄7�����C�6�&��K
�!������qP��nnx-�Gi�1z�!�Y�94��P�ӘJ��PS��Z�Ys!�dÉ{nV)�R��%*U��`�啰cQ��0�Oʅa�K��T@�jZ u�y�"OA�aO�W
EII�6'jtM���'ADb�TD��'NH�*r����R�$U*�T�(���=�IK2I������`P�W�w�:���y�(�ɖ�Z�@'����T�1�VĄȓKj�LB��S�C�䄓�c�� ���ȓ8Lbu��[�9�,{���!׾��ȓAy�%�giV�^y(,rd%$�Be��S�? �l��bO3�j˶� B^�D�"O�i���NƼ�SgE��3$"O�؃0k�pS�@��&H�*̐(�"OH���`��c��A�D�A��'�ў"~�ŃѠL�1�$�1��Id匍�y��B�.�XEY���xC��3�y��T�l�Hxwb�~˖�ٲj��y�F� 9j�� ` 0o����f�L��'Raz"b]	ܒ�C�Cɶx��Q�)\��xR��7Љ�f��4逜 �%�>r2�O���Ĕa"�1�+��P��-	���&�Y��κ8u�u����*	4B��  �����5=���E
|��#>)�4�MË�i�Sn�X��U04$��%�X�!��Ӹ]g�x��NEep���[��Ң%�S�O�` �T.ԿQ�銢m��G˖�
�'$	0p��;euz٨4+R�3T�DP�'0���fDj��#�Ja
�'�:�sǣ�(�q�A,�@�s+%D��Qe�������gء��Õ�!D�8��.�'	�<[�J�e�
�D�<�Ol�O�d�F+҉&W���Ҹ7tm�f"O@��t�ߕmQp�1-Q�l< �T"O���qH
ن!���TO �S�"O��YUIT9Ŕ�Q4�@-���FO�Ujt���� �D/E���2�u�<aq.Q�X��F�L'
)�r�r�<�P��))�e���b��eZ��y�<qr�Z"C���2�Pz��i��Tm�<1g�Қ��`�s��uQ��Bn�_�<كi�:M�j��K&����Y�<y���:F�DI&�ǂwO�"$S�<�2H��i� �dn�;+��}�ugCh�<�Hv��T�"!�����_�<�BH
	fr\� ���>���M�A�<a�E�b���i�,a�Ad{�'7ay���!��A�@��Xv.������yBnR�	��DY��-Q�F�A����y�Co*�H���*���e�3�����<�/Ϸ)�^���N�f�-�%E�X�<��yP�D�񢇶9����ό[�'~ay�+�)�F���l��rb�$)�+�yүA3!wr��w&�2~s���D��1;�����>�$hs(C�H��`x%�`��t�'�h�aW��5�ǥ́[e�8s�'O��(1�ә{�L�F�.Y澼"���d����Q@Ŋ)�H!�j�)�!�D��F�`�q�*�-lS�xa �J�!�D] ��@� ]*;R-ô(X�S�!���ir������q��Ir�Ew�!��5/)�g��\�,�B��21�!�V�(�rVŚ��N��ɋ	h�!���r)>���I?n�V\J���!�Dšm�2p֥�9��X�	�%�Py®����[�{�� �W��*�ybi��;�j!z�)l�z�Ç W �yba	D��a%����ƃ�6���	�D�}�&���t�"]�LX�@B䉾��"bҿJ�0`3p��*4�JC�IjB��c�	<0�
+��@�b�XB�/��9�􀙥y�رr���G�:B�I{�\�Q�S���I0�Ò>o]B��!&�sf�@���Y��S@���D7}nH(}o�D�A%o.,�J�#� ���'�S�π �M��B�\0�}ʳ��sm|	�B��C����G�q6���"(�?�ͺGG�jp��kx� �#F�0&1i�$A4Xqڬ��c�Oآ=�~��O��Q��K4`���ꔮ�Cw���"O2��@nl�Ӧ͜�YG������V�Ou� #k�� �F�RF��H�<��'�����Ŗ9+���`dE.\ ��"�:�"�<E�Dc7xTb�Bt	^�{fd����J�$|!��/#P����u���ړ�L�jf�6O���Ď=lR���J�H��<K�hɹc�!���,<�)���M\��b���(az��O;DO6T���b�����e��!���`
u(Eă@��ux�E^ :؉'~YFy���֛=�d{�BPg�ԺG��y2ț�Q����A�^���G�ɓv��b�Tק��ē2��r��]���ҳ�� ��@�ȓ	uf��b��=V���jB!{�n����O2#<q��4�5b�a�GΉa�l�_����'Ed�HD� |�ҕ92�]�!%n��K� ����S
��D�=z�T�S4�@[������<	���-ƀ0�`�^�qI����h�x�'S�y�ʀ28��	D���k��<r^�d���r�O��������*<��xËT0{�����T�a5��d�Z����7-%*E�u�B�i��v��O�0,I���߹W���FI˔wkb k��c�!�$Ȇ[��yH�N�L�u%%i�'�ўb?�Z��þ�e;�^�	��l` ;D�����[�Z�="3�\({4��Z�/7D���Wg�4%7�Y��ޖ�9J`5D��z�D ��q�	P �\�d8D�t1�.ޯ�Liq�*�=~��F%8��<��G�<T��WLmH��m�<I�J�HbhۃJZ�{`�J��Bi�<�h�.X~�Eh�FG�Ftr�Z��U]�<�drr:�r�m"�q�L�X�<C��Xވ(��ݕH�6�X��W��HOL���ԥ�+2T��a
��>	 r"Ol��3�+p0e����&Z�\����E��~���'w�E��کM�$�,��H�	�'��%��� ���S+0�Գ�}�i����O���q�
����jY���"O��FN�Ca|-���L���A�g NH<ч�R�\�^���aD/c�hijfd�X�'Nў�;�jd8U��b��ڵ���"��m�A(<�s�L�zx>�z�נP��ё	@���'���~
����sJ��bE�
�e���^2:>C�ɥ-��=S��M�%j�AN�,*nc�,G{J|j��M��T%��'�_z�xp��`�� �;;0�h��Xx��;�������ȓ<F�c�O�.�k�ȓ�_�ʹ��3L��B��Q_����LL�������?��ј_���@gѬL��U0�"�D�	�<�QW�HE�4�O5 �$Ż��+R�.�����yb I�
أ�`L+!,ƍ)G�2Q�IA?!�����	�g�5p�Ņ�w�������Ry*B��;T��T�v Z,,�A�a]�Tgh��a؟�������,��Ч͒&'|�`t�/�O>x$�\���Z�хCu�����/D�,Kmܽ�>|(�}΂@&�x�ȓz�����i��^�E��46x0��i$�(1HF5z��[R��.[�����Y&���<c��y�����8�\ه�a�TXHAkML�����ƪ47���:��4��aˆXD��I�	F洆�S�? 2�`��,����G283,y�w"O��7�ΆK(�}Z·'e9E"O��H� B�Ȍ��G�7U�s�"OXp⦯�#ž<"��8��h�f"O½��N�5i2yg�[�v��Q��"Oh}J0���r��8Adخ"��ȱ%"Ota�*�4�8��B3l�� g"O�г@f͏s�|�KVl��|afX�"O�X��Bm���,�K^`0��"Of�r��M8(��d�@�
� %���s"O��JWM��)�&4�7��-L��"O^%��,�0�T���dL1P�L{�<�F,��(Դl���B�-5VmY�Su�<�@��F>D�҇��׾��af�<a "˄y�p����u��r&��^�<Y�i��#E�E�A@�" c���"
t�<�Bo�j
�(��ӚNx���v�<a�C@6��D#$2�ԡ����t�<	�V�]�zy�HR�4oZ|
2(So�<��?/�� �@�����j�<Y�N� %�@<M�h��
�\�<���ؼ����7{~�i9G-IX�<�w�ǕR�� ��.~�&�C�I�<�ᥙ�P�: ��DP�d�������G�<�Ձ@�Sʰ͋pd�O%���A�<���#X�:��c���<����W�|F���h�Z$Q@Ƈ�	� �:���5>�a�ȓ 4F�  �ج�%�H^X챇ȓ�P����E�Ri�a��6X�D�ȓ � ��e���U$� ��<b��ȓH�,��zw4D�#�58[8�ȓC��R�	�K-peK/?�@��#��##i
v�P�V�K%Mr��ȓdv���+zB�T1�!V8G�V̈́ȓ^V���3D�2k1ʉ�G�¶c妴���|8I�
*+Y���wfA-~�Ʌȓs�1c� �h�xz@�é[:p�ȓ\�u:rFE	C��%�>o"��EP ���PA tXBK��n`��ȓk�艉�N�_l}0&�T<[۸��ȓdihܙT��Bu$	��k�n^��8����o��3�L;S��5��JOԼ�w�ʽ-)��H�mƴ7P|��1bvD����FR��C�7	j>��
���Q�t��H�		Jd�ȓr�Ia��ˍ	>�K��¡tpq��h��0Y�eE����&+#[���ȓ�Rd�֮_�*+d���G�B�T�ȓuja��s՘)3լ�5c��ф�G�jA��C�*T�t�"�_�-�F��ȓi��!��(k[���0F_�n��͆� �.A�2C��'a� Z@��ͨ�������@D�XT�Q�"C�m���ȓu:��;U(A�<��8c$��|������#��y|H� aRQ	ZфȓD���w�f���ǭ��U<Fq�ȓ_���P���(_��|S�D�d��ч�78�]�B�D
h�^�B䆐�����s����'x8(�ҩP;��h�ȓb��d���O*�bx��'Ҁ_�H��K������)6��l��RX�ȓLƴ�FN�L����Մ�̘�ٳă�(�0�8���W�̸�ȓ|̔0�`�t�ִ��� 9y�б��S�? @ٹ���Zn��X���
Ԙ�C�"O��۲��*������ۂ���"O��Iᮖ� ܾ�f�A=�84ȥ"O-�1"�\�l: M����0"O~�Q�Ǌ/0<�с�oH(�PY��"On26o�^olm��(Ȕ�Ĥ��"O*8EnL s��a���7"OXy� ��)E�4HƁZ}I��Xu�'\q� c'b�Z�q���4G|,��4ȕ=aW�t�ēs�(4�$80��8Gk�'�"E~Rᑦ;݊Бq���v����$�-B;��j��Ȩ<5!�dU�>f@rd� NLx�k##�D�!��A8�B���)ڧ3�~ ��­Gě3@Z.qք�ʓU��EK�&��mA��2��}Pb�'ي�{%ɗ%��̆�	#'d|�:Dr�ɠ7AF-w���ݱa����e��9T��5�CE�Xp��� ]�44�	�'�>�uHC�v�42��H�N�Q������Y�,(	�A"��O+��"��ϠP=�(�I�M����'x�=£h�q�D�03���STB�2�'�����O�>�9Cj� [ ,��*�}�4I��?D�`C-U�5�S�QF����.}R'��
*�$�M]���w�¹h��fJ�5��zdD,�O93� 	���sa���GT�b��Q�GL@$�jZ��xb	�]H�Y�֩�	��h��N��O��bnB�L7L�>)�ȯ(9a)����zA�-B�!D�P#6�ASE�9 gd��00��cg�<a���D��➢|b��"����	�:PC^�<!�L�<g|K �:#�� '�U�<	q�є@�&����ωMR�Xh1�V�<Q��G;J�@��L��e]~�)$UM�<��b�N���IK�~s�,�1��K�ɖ_��I����׉�ƨ�B�Q2�a��R!��2k�*���8	 ���4��
r�%'���tn��pq��'��!��"�0zdA�5�ٲ{/�Ix�'��5�a��z���b����.}+g�1�Ƒ���n��$քލ-�&�ŬE�9@إ�cE Oj|��\*c%&�J�\#���7`.�{�� �L[F�Q�$D��V�q��*��: �*Y��6?9&)r�}�`�-}��)B����(�m��=ʠ㊤�!�dJ1n�,�s�C)�rh����|�� �N���Do��c>c���A��R�-
�":TJ:�����%a��{Ï��x˦��&b�"�m��F�>5����,Jn��<q���:o��i�Bn-�]q��<O�iÆJw#dx��Lʢe⚼n��E�����3pIdc���C�ɹhvn�"ծ�����!�4R��=�# �Ý*k�4g-N�R�أ|"@�'���a��(*Fn�a��o�<9]-L��9�3	\�`~`y�h��"����m�18��7�,!�y2��L>�M��	��%Iv엪IQ^�)�h�H<Y��ݥi�n$J5F����U[Qk,AD�U�V�#Wi\��!���p=�UcǮL���x��R+mΤ����d�`[VMO�Q�4႑cל�*aB�.�$!T���4C�ɫ4��E��ƿjRQ㢈�?M�8�)Ь��e3~�YUf<K��|"��[#L�RY����CUص��g�<�C��W����Si�_�ʠ��D�4<��!e*;�"t��L�^J@M'?���[
(3e��(Et%���-�O���g��d&�`�Cנvf�}q��)]1�sv���;~R&[6�����W�}Fx��ឧ\���	D�C����S��,���lϐB%H	*�g�5ڶ�,]VBy�̗1/���=D�P�U/1Q�d-�@�"q�&�y�÷>it�\���e)λ���7�8ڧ\e��P���J�F8�	E%:����ȓ$i.I�X�lRģ�Ŕ�7�F�ZJ���7k��Dc���M|�>�%��	2H`��A?r�i�ePh؟"���K���ΊDo&�;!��_��tRt�]�X��B��J�4P;U"O��0S���,��O�E�%�[�q�����"<,b��g�? �����"�fy�K<���"O�:���8�>�H��P�T�.���U��᥉��&�f�:d��.}�R�(<���V�/V��X��ϺsPB�I�)�JD��/U6�s(�RWp���I��
�Ze�;5��� U%'��$��t�r����+g�JY�w�M2�Px�˺L[��ڣ��G����3ɋ42�����<Ny)T*[�:����D=ki�e*��;@4�5K��R���{b���S4ū����ir� Ĩw�y%Gd���D�8D�(�#��g�hC����
"J��7��	r���*�>-̑>EG�F5&r��*�P�:�|T1��6D�<	Ac"6~�L1a�ΎW����O�>�CG���	P��~IzBZ$S��I45��|@s�
��x	�{U�,���pʹ���|V��p����xP'᝹T�����-8�(�b���+�%
���g�џX�+�H�(��9=5��c�9�K4#}p�'Λլ� A"OF�����4hB,)� �P���!�!P�D2�A�b�a�fN����X��(X;�1t��!�-�"���P��C�ɑHG�,�%�W3o�4��2N]���T�O�[0|7͙�sRҁ�S@@~�3�I0<3V����q�����AG��#?���ܽ*�'�����Ī��DWF�tDsJ_�Xټ�1�a�{H���C���аs���"0f��V��~�Ća��!��|1�o�<;�D"��̽N�lpU�Ձ-E ���ۼ�y2-Z��P3��Z+%��8�.����ژ�H�th�w��Ӻ�A�H�Xi/O"�K��� 8���% �1xX�0�'>$QX�!�0{,q����?
 ��*�	B�G�wy���^b�x8G�Q_�'q����� �X[���Pn�Y!��d΂�la������:��0�֨I���!D[U.�R�Nώ5d���� \8la&�3~č���ɠV��'!�X��&��T��5�'�B��rc�p�1���[s,@;��˿�����"OܵT��i+L4�����pb��A���PBo�$���u�>!��^�42J�'Oz�	�mҮ���X���	#{ԙ
�<�� )r�L
RHV�A�F�MV�D��X	)�e�$%���`��TJܱ��c}��[��&�	q�R��Q�J�.]\A!��k�'r���V!���4Y��ED��=�ȓ?~���g�%@�=�.�n�P�ҳX@{�L*���x�Ii���dF0N�@,�N� k]"Q��65�!��'�<�ytlC:n*x���ѥ)�<�X,�D�<����lL����C0�\�0i� 0��R�È�7raz�
��V�D@[?�,���H 0jՊOY"5�#j�&}�qO�� 3�3}�������7)r1�r��&Ϙ'+x-���%JV����O���X���|
`�b�^�#��>) ��w$�U��elE��p?�,ϖ����AX�ڥ�5i��D� ]��M+ k�U����O��� �� [z ���`��<�Q.�/$E��*��)� d��s�<ѲM��K�aá��-1h])��ڷ/ذ���͐�=@)����Tܨi����y�,3jU��<�JB�K'K���$2�7	Wm��,�M������+ֵQ����"<a����20�$�5KW�X��HAB��<9S��Y�l��">q�́�u��9�@�q�H�Ĩw�q�PٴH��u��q�o�y�xg�����mA F�-{%�̿0���C�%�o��dP�DܱR������*j�º#?��߰*���ZqAI�g"��#���=�"��,�; 5�h�+��+���z�w~v�&`�%*��Ų�R�/,LH��'���14��bAXx���kb+�C�6mk��D�@W8��AJ�!���d>OH$8�ł���'���6CG�H�SN��J�Đ�ӓ,����ih\yRem1&��$9Q�qO8b�[�kG^�c�m��Mt� �'q��U>%��E|�gp%ddy��2��(�SJ���2��<�#J[�xt`�Q�B��D{�a3��?����8;�@1Y�Ta2��#�\����c�TAR���dӳk��Y ꂑ#�Tq(&��k�&�VΎ��:<y��`VV���]>��@�#T�Mq�f��<ٲ�^7A��9�F��J��Y!��mh<�f�ܥO���w�H��j
C�Kw�M��`Y*��AP�L#U�8��T'�d�'MDR�%(**2�`ꚏO��Sϓ*):�X��[�I��3e�A�F���"n��|�|<K�o�A�%�$�0�x�� �
�#�@5�F��b߯���N���"�=V<�a�Q�A
l]ˈ�ŭ�D�"!]�V�msե��yҏL�"Ĳ�CQ�^9=d�t�f)XU��8'Ȫ��_;>a���D�փ��O��	9 �mrt�L,z���HRc�&C� C��}�? :��0�߿m,4��q��oQ�P$�C�	u�ݓf"B�za�v��5A#ax�D�E^}�0�B됥����0=	7�H�v�B(�t �!�,8�f�M,F�����V�{��|ɖ'
j��B቎p����Ӄ1��'�H �Rb���'�B�H��]rD01���$�JQ*A��:����3�ǳ%!�$� 
 F9�u�H�BuDP�H�	Yf*�`�T�]��'�����%�<92��)�h��1�^ll�9w�EV�<��#��e�1�X�m�qх���X9��9@l�&�3���\�ay�f
H�V�g��L�i!rk�*۰=Y��Ͽ,@f�r%�/�lp˷
�5|&�i0��<>�s0�&4������T�La���)W���$�:q� U3B��;6���|J��n�P�a�NZy|��Qd�v�<�3f��L�؊��Ahs��𦉒�W	�qO?7�F(p����/�e�\v���%�!�$�Q�&��⩈�es4�D�I��!� �f����G��4ª����E26�!�Ic}R���J$�&�剎�e�!��D;���)�,���ڇ�>�!���>�a��ޭi��m��J�h/!���%h�p�`FYd��W��i!�U�V���o	+\����N×4{!��էW�h��  �H|���-vw!�$� Ld`]�u��2�q�K�-!�ȴm_21��A I�H#Ca;q�!��УiH�`�&:�u�% &.�!�� @``1sDIZ�wH��2 `��Cg!�D�?"��tjR�><xA0D�'Ex!��;#IԑI�
O*!?P��M%4�!��'i�n@����A.�#�ѩ6v!�$Sz֤���G1�,�K%�!� �H<��i�䅂���GH΄b�!��T���a0	z� �ٲ`"!�$�Q"D]���c�|�Y6�[p�!���dwTz��-��"��ڛU�!�d�2�re
�( ��5���Vs!��8ISڐ:��ޫ9��Q��bS!�$R8 �lIa\ b�X�c#o�2$d!�B { �IS�g����׃>!��פ3(��w'ոLt�I*6kM�!�]���� ܰ>ٜ|�"GD& �!��= ��I1aG��Q���Y��!���#g��Yg�N�V��(zAhK�f�!��o�8	�&��PqB�L�<�!��9����#�G�E�j�(���
zy!�D�*wJ�9�ܰ3��4k�G��r�!���tRua��Y�p`b�%�X�!��=q�� ���1�`��d�&�!��d�xP�@�L���04Û	�!���W����/@�n�#� -�!���
a��R!�}���
D �!�$�<;VP��sB��p��iۼf�!�$@�S�4�0�S8J���5Ɵ�!��S�f`ʡᣣ�W���I��D�[d!��НB؂(�AA�&�pp0��߷oi!�d�6�V�K��:E��l�ԍD'VV!��\>����բ��xa��2dN�8Lf!��ʛT �� ?"�l�)Q�R�3!�$�-����4h�&gz9��̎k!�D�'08�Xs%�9ndI��D66�!�M�i��8� cA�Y�����
��!�ę5�X}�e.� %yp`�.�6)Z!�Ĝ>"� *�~65�WJ�$0!�$Q�e���IՄ�GB]�qd�,
8!������#צ'h�x����(D-!�� ����ӮX��x ���6	ؤ@q"O��qd�4F=p��/��.����a"O�E�#㑢���� /��R�0�0"O&Ex̈́(��]s���=a�`kT"O�5�%�BHz C1M�1Dn�""O��qv�²�+��?Y60��"O�	iq�Ӎg��(r����^C:EW"O�ը�*����&A��R;d���"O�4��|��\h��ހ�����"OVy�tk����Jd�MCvTj@"O��h��/VK��-E�RD�H�F"O"A���׉Y�
���.R��0r�'�&I��`��3���N<9���
�O_�P���ē>S�zjEXy��BE(o�8LF~���R.��ڃ�i�(^���' ���l�:�!�Ăf�����
,����2ʉy:�D�?Qn}�dF���)�'a�=�e�S�)����N2$oZ�� 8^��g��r�%�F1����O��{bA��g.�)	Ó4������':���#/Wc{����I�1�Ժ�T>4���I���>L8<����<AbX�k#OĲ�O�/w���i^8c<b��!�ɬI'�d��g�9�1������a`���6��)��"O:�� /��Kxp���
� #�U���O�H�#�E>*ZnI��}:�A'�|J��Q]/�� *U�<����Su�E0]P�ht�L��N�5h���Q(�<�0<A��Þ �b�S�����D�E��$A!���|���&�&o���;�.Yj����lC!�$�4}��8�e+�,��˕a�3V����{deA�Yb��}��iI�M�X�C�IŘ\1T- ��r�<	�����eY�>*;���MMKy�%������=E��H�J<�E�.&>1������y���V��
"c}jؘR��1�yR
�e�����_�\R}��,��y��PnP|��@ ��W�`��!�߰�yr���`�Rd� ݐI����̈́���!�t��7B;�)����Js���!��D� _�B�	�/�T-��G܈L� Ů] 9��J>�.�;�>�OnI�7%	.:|ū���Xʴ��OlA�W�T�O&��T�O�`��k�kΧ�B	�$���p?��أ)�lh�H�g��:Qc�_�DQC��CJb%k�>��A�:7�^!���)S����r��U�<)�/�3_j�Q Ġa�(�4�Q~�$��D	���ɒO��'S�t5���R"c����nZ;*�,C�ɀ0�FhK$#�24�\Q��B�I� S�>�&�4%��!�|�<�4��?]hF��d��RK��sç�b<�dL=0}��Jqd$Y �Ȕ�6_#�`�^-B�H��A�	��=)SF�.\�{d��<(�y!y�� Y!.Z$�a�M[)
���!�4/���1E-���#�3,����6hd��ɐ	Y���(8�p��'4"�FU�Ru8���Ì[�1E���	�gt1)���Drpu��y2G��w�P�8�T�S^X-@��pq|;7KD�G�@�nZ��*$V��|�%B�" �iв˚�B��d@����x���4u ^��휟]�,�Xb���q�JDC'�ՋL��ɹ��C
'��zh�;:Ӳ&H:�z���l��0>����bt$�0d�� ��ɡ�Ń1*�칠s���:�.݆�{�t!��	IN���j{�y�'��b�cC<~��(��/�0G�$�D��j� ��Ё7��� Ī(�����y�n*�N8��Mƿ�<�4���Hw��X-��f��U$@k�M�J�3�ɻQ[�Ē�W ?�I�1.�2X
,��du��x����-���N�V��P��нK�����!Qo�|B�O0\O���� Oظ���ã''TS��dOX�1c
���P �Q���ʜΠ�#�J��KR�ЊVs!�$�7r,���
o(LDԏds���W��H#�bS!|�0$��-
8��>��E��@W2$����~ �1���.D�� ���'.��c��,yB 	.�̡��$8}҄DPJ��/)��D�Q��`��� � a��׿oOa�MI-�z�����7����@ ;�U��$B���I-����)�	�
X������"?q� �K�h������6��!(�+P(h�����-��� l�v"O�ؐE����L!�吥%L4���Q�5ʙ�.� 9q����gfزT�k6,��F��h��s�&�*G-,C䉳|Y���HK�o#fh�U�s��0��PM��\�6B6Y���wO.�� QX��R`Q	� ���|!�$�S����лV'.|�AL�;.<��UIܫ3 �+բC��|1�����rd_�GE:�pqh��~����C��~Y��̐�MSP�C35�D��'d�1�D�:��t�<ɴ(����ڃ$�]!���r@Nh��V^ �ie�ж&�#}�� "sb<��D�f<����*]Q�<9��Q7V�i]: h�� w�ټmq�#�H���h��P�Zv����Ѭ���c@;_]!�$А[t&�f��\�C�-E�&)�|�$%¡i���Q�D9`�Z���	ly��k"U��è��'�n;��2�ȕrj��?r��7J����硗'5��A0-E~��B��
BU'��!���S<�8S&,01��
z�±@G���"~�q��Gi.e:`�����-v�=D��)��N+5Z5�ŎӪ;?��6+R�B��q��aj���<�j'>c��#�h  ���CAQ�8l�� �D��TL0}�"@=�p�vD >r֔U��.8PVC�h@��I)Q-f�m�P�h�a�P.e��	�i���BMC~��ֱk�(yQ�.Z�S�� ��g/�>,�\��$R"QL`C�	�Lwڭ�@ɓiؼ�C�,\�4�K��h#`�L!j�,O��	4jМ�A�<Q���3������h�4��J��t�$b�9� E���L�7 L�ȧ
-_�֍X��C�I	�	*r�l��b�'Wџx����>�hx'<f΁��.*�.7� ���ʓtS��h���=����D��
��-�@l�}�>����<�ON�H1N��X��^�#/t]�?O�\ɀ��g��*�O����^�`�pc>���e"IR��Rã�1A�Z� �3D�4(U��=���r��?I���/?ɕ���� jZ�'�֜2'��E�$C�i��XOW-8���@�O�a~�'f�eC�bs6��_�`h3��i-.(���ɚ�@&	��m�ǗhH�\�>��e��1�Zp�G�V�z�.���i�wD�#�
]�u� A3� �y��ۆ(0�ܹ�A��vB��y0��b��y�"�I�Y��J��O����Y�PB'E�V<�`�	�%L�}���9D�t�A%�('0�M��e�t�P%�`�Q�JrC�YR�P�Mrx���dMٺ|��yX�"?N���5LO8�:a�ϓ/�`��'9���5*�jٱ�)B�����=�� WFt��OR)1��;#Ya�#H�\`���dDP�B���~b��;C>0�O�h�P�T��Q��j͠V8^k �!�Ӫ�p?�FKs���e��}�F�Ae	i�LI)a�m�l���ԜW�J��'9m��
w�S�o�t�n���Ǣޟ(=r)���\��`�h8D�,8���2`D�����ת� �cք�ɘc�$
�\9t�.Z�1s�,� fΌ�ɮ�:&`�2%��DO�j)V�n[�r���hv U�az�-�8JDL{�*�Ɵ\k���-�A�T	ȭJ�h�_K���!��N���1s �e��N/��O��wm�9�dE���0\4���v󤂰^2���'��?�Q�ֶ]�0(�Cl>��mͷ⨽��.�^�I "[�R�L���
3Za~�,� `�Q��D���b�	�,t�H�zQ b�`�+���F�J�<�$t��I�B���r�),�y��rY��ϋ�9�pʐ"�yR��< s�� á<o�"�͍�R���;0݀4�s������u'O@�<�'B����:O�Ä�\�f�ʑ�F-U�ErO4�R$#�&�6���6���w�"E?­9¯���y��+s�.4b�c�Z�'��	�kO�%5\RU��EEv���I`4��J@1���	�2t
�)s���5p�'�١�Kxh[�\xp�����^���#".�\5pM&��3b�C+^1tI�'�~�B��x�S$qHR��ê_:fy�QK�e��C��"Zh���J�m� y�0f\��f%���ʂg�>�]llMC�m9X.@�sK;Sg�\�ȓK"��B��Q�Ȣ��ݰ$�9��S�? re
�ɒ,*���sK�$�y�5"O@��"c�
'�~�K JD�Os��c�"O��{�E��1�j�Y4���!�"O촠��URKԁ�dF@�y��@"ON���NNM�v1���3o{DhA�"OL=�M<[�~ӏɁD3|��"Oz�!��E��d�qn�=+��!�"O��	 !��}��ҔL4v>���"O�����֑z&1⒋T.��9�&"O|z�̑:NS<lr�)ӓ{�
&"O��s���Q���9N]u�d)�"O�!����'T����,tRfh�G"Oʬ0�Ɲ�,��D u�߲|?��3T"O�p�ïŲ-,D�B'�ەs,t�K�"O�E�F�@�g�*\9H��cz�-hs"Oui���T�C[Z_�Ͳt"O��cDE!�D��-; L� �"O�89D��,�A�c���p#ެ�w"O�����VJ�*������G�t�B"O8���w�6	+dc95�^�	�"O(5��M��}ՎL��]�Nn�h�b"OP����#Vz��Q� TJ�B "Oph���P��!��k9P��"O<��Q�ۻ{:*dbF��
\�}�<�v�� �T(&��{�2���A�<��C�>v��Ï�P��Ȱei�~�<���=iy�1���Q�Z��07	[y�<�ҌJ�	X����ם�D\ 2�@p�<)F)��^���poPg��{�N�H�<���}�~� ��@��öIR\�<�sǙ�f��H3��I�\�Dd���NR�<�qaV��-)eKK�P�P{uJ
w�<�B��-"�l�Tg�6,�^xX�_�<��a�e����D.O����_ک*�k]=L���.a~]`��8ڧ73r�싓�t@���4�BEq#: ��ʓ2���OW��*�B�NF�s`��^�Tђd�iyb���3	x%ZUk2���S��F�NxՑ�ϝI�x�h�W� xҋ�,~�6L�֣��0|a�I�V�`��#��u(;�CEަ5aǪ�lSx@f�Ney��	U! Ø�fB5tG��!5̝�<xR
"�^h$PK/O���Ӡ`N��i#�?l�r`Id�=Z����I6���Z�jY��'s����H[F��\+#H}9�(�<�gT�p��(���t��'۬Ɉw�I1Z%�]�#-ͶM��QP�OH��2gm���O>ݲ� �T�0�X*��Ԝ!3�׭�M��JZjB����Z?E�TFP/[����	�M��Y�F��>��ȱ�e�+��h�+�h%��(̜+\T���ӓk�l��jB�84�穟9A�9��;*�$�A��|����0�<�i�@/K2�ye��Xf�6.
�4ØW7UI� eWa�d��$o��u(𢞴�8�2ҫ�-":L��
/�M�A��#���*
�'DL
�'�ڱ �9SY�o!0�HԄ �qS���:}���iF���.n_zT��ˬb^�Pjp�͎ R�&�\m:���'�������Ի�BL��j�����M!j>���ĠT��P[�k���.��f�1?���2�Y���,��)CO�H�A���=+D)�̡Da�I�7��Q1j�o~��Z�I52�K>}�i�RM@	�%���V�!b�p���6(���'�p"}��O�N< ��(G��೐`,gn@�$ʄ� PH�zD
J�<�b�F�0|��ܹ��f�xK��Ch ¤i��ݛx EhF�7$�<���{�d��8ι����9`�D�W�
�1�l5����+����~B��)B/���B�"U�_�4+ �X� �R�\�D,PA�J3Ӓ����l��x �7{�%�E�O�n�by�v�=Q�&����c��R˳|J��͊e��R4��;!�rP"�o�G�<��L:88���2{\Jd2WM�<��[�8���$-��'�j�ɳ�XL�<�1;���s��*n̈́l�p��B�<)E�:P�X����
��$�}�<A��A5Ⰲ�Ε#�"��.�z�<� ̐:�GL�o�.�2w��1A�"OB��vc��6V ����[6i,�g"O�Yk��A�IȂ�#�J	Q��T"O���o�����Z7��[p\�"O���5Ƒ�+�R��7ɗ b��QY�"O<��$�D�^:�|�3(W��HK5"O�(���h1�M�t&נJ�Z���"O�L�c�,ST jre��5���	a"Or��JU�8��i�����"O,х�X�fybȳե�?h~TQ�D"Oh��&�#b[�R�MV�$��"O����+*�t;��G�x�<���"O�U#��\Ҟ�
�	BoXl�4"O���B�[]�u��Ol��P"O�AI!��_w$����9h5  "O��*�/�¹Y&@�"��2"O�@�u�B�s�.4����vH;�"O&(9ר�)�̈
7�פ!���"O�xp�Bˀm�����-<��3"O6Xx�q�� eDʃC$h��"O2�qP'�/PU�% ��$�ErS"O�I���P�"��acۉ�J��V"Oq�G�4:�: �,��k�� !�"OXt��	�hቇk�(
rՙ�"O��wҾ"8L(��CѣY��0"O��i"&� �`	����%q���q�"O p���G�xJcaߔ1�d"O�ݓ��.cݐ�@ �	Dφ��"Od\S6JH,"�rL�5EɀB�rY��"Or�:u�0?���S�j�61ވ5��"O�	� 쉻�P��3�1#�n-(�"O�Q2��^f�ք$��2H��(4"OV��� �.Q1�ϚA�!�b"Ob�Q��,�S(� Z,��Y"O���q�E0S��-�gF�W(���Q"Ozm��c��<R�E��j� �"O`�J@k����`Re�7�3r"O*�p��4qC¨�c�� ,��Q��"O�����B18l��o�*��hr"Opy8c�S�Z�ڠqu��6�.�4"O�d�(�:�,�JGiY�'器±"Od�����xbt�
F�X�q�"Oj���HF;rvQ�����<�� �g"O S��ٱy�c�����s�"O�X���K�4�"@$^
,;2�G"Oz)����|�� �� �"Ot���]S�ν�P���*�૴"O���
Ы%Y�`a L"x϶�:6"O�A�&�|�p�$�ц-���c�"Od�xc�̖k
�u3F%��P.���"O�:�M u�����+
����"O�H�F�JT�M;���4�)Q"O0yQd+�Lq����I�X��8��"O�D�Ӎ]�(�ЛS��)>��"O��[1��0��\���H-'랝*7"O�Mc@��-��|C& 	7W�=� "O �C��{I@ۢ�$O�
��"O,�b�oV�*?4��U
Z�,�� "OL�u��x��lH�pp��x�"O~�9�/�xg ���d�;AL=�C"Of%B�MP.n�!�A��S��k�"O�$�qˇ)�\	c��6B����!"O�XbE ���: c��A�P��,	 "O.��w�W>e�P��R�J0z�ڬÁ"O� �$ �c�3�%�A*�N:�;�"O�1SE �3�����B�>l��"Oz0J��Qv�9��]��tS�"O��zp��5/~ZlU�!�JhQ�"O&M�ϙ� ��AAL(#���f"O8�E
�:$��ёŞ���XD"Oxc�&T�oC��M�/�i"�"O��R��&-rZ<��l�!`^2Lx�"Ob sd�B��!�b�rcNسf"O~)��N :і��#!M�^NIp"O�Ik�	لmca��}A�q@�"Oh���,0��@w �8R�h�'"O��iDk��)D��С�\18c�\˓"O��Cs�
8��	��ڤ�N��"OZ�r���h2���� �|�"O*q�g�0{Y�$)��(H�0x�d"O|y�qlٯ����&�:9�J�C�"O���bޡ#��`S�X��,�"O�i+���O��m���%n�R,�u"O��3�$թg����%�H!oϰER�"O��˧���8�>�HP��"O�U23�R�ND�Y!��%OW�yBA�,."hхKD�zY����OA��y�*G�=+�h1�
�a%:�Ӧ��yaΎy���ď�2j2��E�y"@լ#�l�s���LP�b��<�y�I��=�2��ض{(�����yr�
�F	J�b�� p�q� -�y��J(�a�����X��aԞ�y"NWJ�90�ģPD!c!D.�yrl�	�hr�� \4���dͰ�y�B\)Q\2�a�MK �! Ƈ�y�ᄕP��L��*�x)�4���yR��1"����i�	�*9�G�] �yd(:���o�nm�`ȷ����y��R.�Ft�ed�!�0���� �y�B�`��a��1�~�H����y�A�
�t$��!B6��jrh�y���2�����M�0 ��	�0��y���/�������pi�Ï%�yR�كA��I��AR��lY$B
�y�I\� R�Y�IH�R��ƒ�y��A�z�rAV��ҭ�����y�f,̰�s�a�{���&M�yRn�$ u�P�lýsd�ຢ�͌�yr��L�
U�6�8�
�>�yr	Z�D����؉%����f���y�N�9J�&E���S�$� �e����yb���J,���e�^�q-R�`��	t�<9���.,A��1��4|X����c�<�P蓜)vq[�b�z0���^�<a��EM�4���Μ-��-�A#�C�<9G�1 #��aCu��%.A�<q�h� �!��$�}�dd�F�MB�<1R��-v*�c6N�I@شC�I{�<I�.I�s��A�S�	��Ě�@�r�<�ub@�7N�)�;18����v�<��F��M�5L1w�Jq���n�<�I$ �����!g��X� CC�<��%I��ƤHX��l��J�<��Aԍ)�*����6Y�G z�<Ya#��X"�pI�X�:q���v�<ٱ��,{�K�o����lRDK�s�<����nXv�#���5��l�<� P )�?�>�h�@%@v�S�"OJ���(D�y6,9$'�.�n���"O%@e$�txm�@e�
�`y�F"O�0v���r�4�r��_�|sP"O�	s,�!A�3 �Z�;"OP����7�\��!ޫ3^���'�<͂��
_kd�աO�fV�H�'N�2��ؼ)�(�q���N�����'M����Ұ�8i��t�4���'�T��Ο�"q�����R�:P�%��'�+$�!W��r%hHE���'���L<%�2��sL�9RT`�'�BT
a�L�9�gP10����'e4�����p:Ҹ!��¬;yZ\��'
����K�
�����Q�-��ݰ�'o@0�G��5]������P���y�'��!�rǎ�/S �����E5�I��'b�� �2 ��@�hR�9&��K
�'����7�������Kc��	�'�8]!�� 8�Ԑi�]U���	�'�p��ŋ�VϨ1P�J(�4M�	�'��D)k�6wn�r��'����	�'[�b�B�mBL�:� ���K�'�Rͣ��S<*�8����-<�f�	�'<��s���)�t�ҵ�Q�-,Y��'-\��7!�Y$��S�M
*\����'��MJ�`Q�|@��Se� 4|X�'��ss,�
.����%��$���'1x��#L�3���k��K�kp�l��'N���
,\��(F�	q:6���'o�k4b�*���)%�O-y� ���'��!%m@�~����N˂l�hܑ�'}����@_qk�	�7��0�Bk�'�`�zEQ�,X�. -��}h�'�b|pfh]{���"#�ɑ�'�na(Ц�)POl�ҥC�	�'�VE����x["``6O�f�8���'ܾ�3%���+3.��̛0~DtI�'������R�Su �T�ݦV*E��'�$�%�ͬb��Db�ច!�k�'�4A����� D�ĳ�$Y�'�(dفBٝ�xM�F�Z
վ�b�'�Rd�w��o�5�W3�����'*]���Ô2�ҩ9Sc�U"���':�,�0%<Z ˲��I�����';���f�?���bK�/2�$��'��`�6g
�ex���k�*W�h��'���Ǭ߃t���D�V&RX�8
�'��	����(���K���	�'���bq����v�A?��T��'9�y�Y:RLT!�m�,��
�'G�|���*n��� ��٢j-����'}�D�#��/�&l���_�^yX�'Қ�{׌�91[�|su�(Q.�i�'�6P�M@�
�l����^�x��ܣ�'_h�!B�7��X@V�Vb�(�
�''������!~V	��.�^M)
�'ĜHD
.3N�yp����ڼ 	�'���8�jEMd�x��݊N�y�'���Z���?�9���>"�py�
�'��(h�a�16�u;5˘� � Q�'*4aD̒H��Z#���0�
�'��'Ц+x(��^&Q�8V��>i�18\��-�q����Z����v��0d@"��p�4��/T4Z�=x�"�>DX014ޟh������� �Ŋ����c~�ij5%B/r��:A(ӰB@8���<BT��Z%��(��O�t��FLJcL��I*2���0T)��i�%3Ǫ\�N{t���Or1JF�'�J?���O&��n���U�I-W1��J�|2�m
��>��nrz=s@;CԸLz�mH?c��e�� ś��'�ɧ�T�'���4y��A7�bD�Q�_p��$+Z �M���?qlZ(r��D��d��PL�l���A�J4ʈ��N^n.�p!fA;z0���e!�U���r ��%��uZ���>[�Œ�8P,��Ѿem�\�Rc5y�9J�ϗڱO�H���i��\�ÆWk�r4�b�Z�8I:�Ei�)l�%�x���?�'��'9����K!j� e�HPai�'��1ۥ�ǣO� �X���5�����������M���?�'.}����P���'��Qac#h�������P\��$�O�h@eWh����oM�'Ӛ����7@$��͌�s��EϿ؂ђ��D�_�{��Խ�Q�
؊IL���J@�E�x]��¢JU���t$Q'���7
�L�6�ā��ҟ�r�4�?y^w��s1��!���bs�v>.<��'����?�'��C
U�z�%�W�a��e�D�6�O��lZ�R��$���߃����A�Q;3�^�!
oyb�T!Z��6�O ���|b�!�+�?��4
�C3�Zo|�]��� ��`"q�'Ra���\Q�0�"��&���#�E�,��֝N �"��Z�*���ʀPͮ�8�O��a q8�c���;?Pn "քX�"9�1R��,�č�$"p��c%��h�>x��P�����+���'V���b?%ٕ��9;.(l��(S�w�l��w�&}�'�a{2��Ul8ms7��5{�B��rM	�~2�DΘ'�@6m�O�b?��fS�X��K�B�	�Pi`�/>�?1,O�����	E~���-�(��5��m��E*�����JPrqNi�|���.Q�N,���O�tm�m�kc-k��$6{�9#!������� ݺd��+Pa�3,�!iF�#^KX<2�b�F?1�֑O��LT����h4xRc�:S�t7��OX:�o�OFMKO|�'��D�i�p@���B�[���'�
(y%�(��'a"̛~@�1ciR5n����k�����hӶ�D�OV�l�X�$�'��S6��󀚠i4NpPb�Q/iЊ��F�M��џ|��ڟ�������O�<P�N��zqXE��p���{AIYo�0�;�MٜL5�=k�Hң�FI���d�X�.��㫛"l�fi�co1
(:`�8>�0�k��ۜB�E��%μ�z���?�	/@07MZ�e��� &-�`uz'�D=w[����-�M�����$�O\��I��	�ա2z�bd�)@BqOZ�=%?Q˂#�$W��S�&��rm4��`)}r�j� ���<����?	����M�w� �  �